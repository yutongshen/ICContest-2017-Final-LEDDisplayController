
module DataReceiver_DW01_inc_0 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;

  wire   [9:2] carry;

  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[9]), .B(A[9]), .Y(SUM[9]) );
  CLKINVX1 U2 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module DataReceiver ( DCK, DAI, DEN, rst, addr, data, en1, en2 );
  output [8:0] addr;
  output [15:0] data;
  input DCK, DAI, DEN, rst;
  output en1, en2;
  wire   in_cs_1_, wd_addr_9_, r_data_16_, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, N34, N35, N36, n1, n3, n6, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n350, n360, n37, n38, n39, n40, n41, n42, n43, n44, n46,
         n47, n48, n330, n340, n45, n49;

  DFFQX1 en1_reg ( .D(N35), .CK(DCK), .Q(en1) );
  DFFQX1 en2_reg ( .D(N36), .CK(DCK), .Q(en2) );
  DFFRX1 r_data_reg_14_ ( .D(data[15]), .CK(DCK), .RN(n49), .Q(data[14]) );
  DFFRX1 r_data_reg_13_ ( .D(data[14]), .CK(DCK), .RN(n49), .Q(data[13]) );
  DFFRX1 r_data_reg_12_ ( .D(data[13]), .CK(DCK), .RN(n49), .Q(data[12]) );
  DFFRX1 r_data_reg_11_ ( .D(data[12]), .CK(DCK), .RN(n49), .Q(data[11]) );
  DFFRX1 r_data_reg_10_ ( .D(data[11]), .CK(DCK), .RN(n49), .Q(data[10]) );
  DFFRX1 r_data_reg_9_ ( .D(data[10]), .CK(DCK), .RN(n49), .Q(data[9]) );
  DFFRX1 r_data_reg_8_ ( .D(data[9]), .CK(DCK), .RN(n49), .Q(data[8]) );
  DFFRX1 r_data_reg_7_ ( .D(data[8]), .CK(DCK), .RN(n49), .Q(data[7]) );
  DFFRX1 r_data_reg_6_ ( .D(data[7]), .CK(DCK), .RN(n49), .Q(data[6]) );
  DFFRX1 r_data_reg_5_ ( .D(data[6]), .CK(DCK), .RN(n49), .Q(data[5]) );
  DFFRX1 r_data_reg_4_ ( .D(data[5]), .CK(DCK), .RN(n49), .Q(data[4]) );
  DFFRX1 r_data_reg_3_ ( .D(data[4]), .CK(DCK), .RN(n49), .Q(data[3]) );
  DFFRX1 r_data_reg_2_ ( .D(data[3]), .CK(DCK), .RN(n49), .Q(data[2]) );
  DFFRX1 r_data_reg_1_ ( .D(data[2]), .CK(DCK), .RN(n49), .Q(data[1]) );
  DFFRX1 r_data_reg_0_ ( .D(data[1]), .CK(DCK), .RN(n49), .Q(data[0]) );
  DFFRX1 r_data_reg_16_ ( .D(DAI), .CK(DCK), .RN(n49), .Q(r_data_16_) );
  DFFRX1 in_cs_reg_1_ ( .D(n47), .CK(DCK), .RN(n49), .Q(in_cs_1_) );
  DFFRX1 wd_addr_reg_9_ ( .D(n350), .CK(DCK), .RN(n49), .Q(wd_addr_9_) );
  INVX3 U4 ( .A(n1), .Y(n45) );
  AOI211X1 U6 ( .A0(n46), .A1(DEN), .B0(n6), .C0(n45), .Y(n3) );
  NOR3X1 U7 ( .A(in_cs_1_), .B(n46), .C(DEN), .Y(n6) );
  NAND2X1 U8 ( .A(n46), .B(in_cs_1_), .Y(n1) );
  OAI32X1 U9 ( .A0(n330), .A1(in_cs_1_), .A2(n3), .B0(n46), .B1(n340), .Y(n48)
         );
  CLKINVX1 U10 ( .A(n3), .Y(n340) );
  OAI2BB2XL U11 ( .B0(n46), .B1(n3), .A0N(in_cs_1_), .A1N(n3), .Y(n47) );
  OAI2BB2XL U12 ( .B0(n45), .B1(n8), .A0N(N33), .A1N(n45), .Y(n360) );
  OAI2BB2XL U13 ( .B0(n45), .B1(n9), .A0N(N32), .A1N(n45), .Y(n37) );
  AO22X1 U14 ( .A0(n1), .A1(wd_addr_9_), .B0(N34), .B1(n45), .Y(n350) );
  OAI2BB2XL U15 ( .B0(n45), .B1(n10), .A0N(N31), .A1N(n45), .Y(n38) );
  OAI2BB2XL U16 ( .B0(n45), .B1(n11), .A0N(N30), .A1N(n45), .Y(n39) );
  OAI2BB2XL U17 ( .B0(n45), .B1(n12), .A0N(N29), .A1N(n45), .Y(n40) );
  OAI2BB2XL U18 ( .B0(n45), .B1(n13), .A0N(N28), .A1N(n45), .Y(n41) );
  OAI2BB2XL U19 ( .B0(n45), .B1(n14), .A0N(N27), .A1N(n45), .Y(n42) );
  OAI2BB2XL U20 ( .B0(n45), .B1(n15), .A0N(N26), .A1N(n45), .Y(n43) );
  OAI2BB2XL U21 ( .B0(n45), .B1(n16), .A0N(N25), .A1N(n45), .Y(n44) );
  NAND2X1 U22 ( .A(n6), .B(wd_addr_9_), .Y(N36) );
  NAND2BX1 U23 ( .AN(wd_addr_9_), .B(n6), .Y(N35) );
  DataReceiver_DW01_inc_0 add_73 ( .A({wd_addr_9_, addr}), .SUM({N34, N33, N32, 
        N31, N30, N29, N28, N27, N26, N25}) );
  DFFRX1 wd_addr_reg_2_ ( .D(n42), .CK(DCK), .RN(n49), .Q(addr[2]), .QN(n14)
         );
  DFFRX1 wd_addr_reg_1_ ( .D(n43), .CK(DCK), .RN(n49), .Q(addr[1]), .QN(n15)
         );
  DFFRX1 wd_addr_reg_0_ ( .D(n44), .CK(DCK), .RN(n49), .Q(addr[0]), .QN(n16)
         );
  DFFRX1 wd_addr_reg_3_ ( .D(n41), .CK(DCK), .RN(n49), .Q(addr[3]), .QN(n13)
         );
  DFFRX1 wd_addr_reg_4_ ( .D(n40), .CK(DCK), .RN(n49), .Q(addr[4]), .QN(n12)
         );
  DFFRX1 wd_addr_reg_5_ ( .D(n39), .CK(DCK), .RN(n49), .Q(addr[5]), .QN(n11)
         );
  DFFRX1 in_cs_reg_0_ ( .D(n48), .CK(DCK), .RN(n49), .Q(n330), .QN(n46) );
  DFFRX1 wd_addr_reg_6_ ( .D(n38), .CK(DCK), .RN(n49), .Q(addr[6]), .QN(n10)
         );
  DFFRX1 wd_addr_reg_7_ ( .D(n37), .CK(DCK), .RN(n49), .Q(addr[7]), .QN(n9) );
  DFFRX1 wd_addr_reg_8_ ( .D(n360), .CK(DCK), .RN(n49), .Q(addr[8]), .QN(n8)
         );
  DFFSRXL r_data_reg_15_ ( .D(r_data_16_), .CK(DCK), .SN(1'b1), .RN(n49), .Q(
        data[15]) );
  INVX6 U3 ( .A(rst), .Y(n49) );
endmodule


module PWMConvert_DW01_inc_0 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [16:2] carry;

  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(n3), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_13 ( .A(A[13]), .B(n4), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  CMPR22X4 U1_1_7 ( .A(A[7]), .B(n5), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(A[1]), .B(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDHX4 U1_1_9 ( .A(A[9]), .B(n2), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  CMPR22X2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX2 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  BUFX8 U1 ( .A(A[0]), .Y(n1) );
  INVXL U2 ( .A(n1), .Y(SUM[0]) );
  AND2X2 U3 ( .A(A[8]), .B(carry[8]), .Y(n2) );
  AND2X2 U4 ( .A(A[2]), .B(carry[2]), .Y(n3) );
  AND2X2 U5 ( .A(A[12]), .B(carry[12]), .Y(n4) );
  AND2X2 U6 ( .A(A[6]), .B(carry[6]), .Y(n5) );
  XOR2XL U7 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XOR2XL U8 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XOR2XL U9 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X4 U10 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  XOR2XL U11 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
endmodule


module PWMConvert_DW01_inc_1 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;
  wire   [16:2] carry;

  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_1 ( .A(A[1]), .B(n1), .CO(carry[2]), .S(SUM[1]) );
  BUFX4 U1 ( .A(A[0]), .Y(n1) );
  XOR2X1 U2 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2X2 U3 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  NAND2X2 U4 ( .A(n15), .B(A[16]), .Y(n19) );
  NAND2X6 U5 ( .A(A[15]), .B(carry[15]), .Y(n15) );
  NAND2X2 U6 ( .A(carry[16]), .B(n17), .Y(n18) );
  INVX1 U7 ( .A(n15), .Y(carry[16]) );
  NAND2X2 U8 ( .A(n18), .B(n19), .Y(SUM[16]) );
  INVX8 U9 ( .A(n10), .Y(carry[6]) );
  NAND2X6 U10 ( .A(A[5]), .B(n7), .Y(n10) );
  INVX4 U11 ( .A(n16), .Y(carry[14]) );
  AND2X2 U12 ( .A(A[4]), .B(n14), .Y(n7) );
  AND2X2 U13 ( .A(carry[8]), .B(n6), .Y(n9) );
  AND2X2 U14 ( .A(A[2]), .B(carry[2]), .Y(n11) );
  AND2X2 U15 ( .A(A[3]), .B(n11), .Y(n14) );
  AND2X2 U16 ( .A(A[8]), .B(carry[8]), .Y(n2) );
  AND2X2 U17 ( .A(A[8]), .B(n9), .Y(n3) );
  AND2X2 U18 ( .A(A[11]), .B(n3), .Y(n4) );
  AND2X2 U19 ( .A(A[12]), .B(n4), .Y(n5) );
  AND2X2 U20 ( .A(A[9]), .B(A[10]), .Y(n6) );
  INVXL U21 ( .A(n1), .Y(SUM[0]) );
  INVX8 U22 ( .A(n8), .Y(carry[15]) );
  NAND2X8 U23 ( .A(A[14]), .B(carry[14]), .Y(n8) );
  XOR2XL U24 ( .A(A[5]), .B(n7), .Y(SUM[5]) );
  NAND2X8 U25 ( .A(A[6]), .B(carry[6]), .Y(n12) );
  XOR2X1 U26 ( .A(A[10]), .B(n13), .Y(SUM[10]) );
  AND2X2 U27 ( .A(A[9]), .B(n2), .Y(n13) );
  XOR2XL U28 ( .A(A[11]), .B(n3), .Y(SUM[11]) );
  XOR2XL U29 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  INVX8 U30 ( .A(n12), .Y(carry[7]) );
  NAND2X2 U31 ( .A(A[13]), .B(n5), .Y(n16) );
  XOR2XL U32 ( .A(A[3]), .B(n11), .Y(SUM[3]) );
  XOR2XL U33 ( .A(A[4]), .B(n14), .Y(SUM[4]) );
  XOR2XL U34 ( .A(A[12]), .B(n4), .Y(SUM[12]) );
  XOR2XL U35 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U36 ( .A(A[9]), .B(n2), .Y(SUM[9]) );
  XOR2XL U37 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  CLKINVX1 U38 ( .A(A[16]), .Y(n17) );
  XOR2XL U39 ( .A(A[13]), .B(n5), .Y(SUM[13]) );
endmodule


module PWMConvert_DW01_inc_2 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [16:2] carry;

  ADDHX1 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(n2), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(n3), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHX4 U1_1_1 ( .A(n1), .B(n4), .CO(carry[2]), .S(SUM[1]) );
  BUFX4 U1 ( .A(A[1]), .Y(n1) );
  NAND2X4 U2 ( .A(A[2]), .B(carry[2]), .Y(n5) );
  BUFX4 U3 ( .A(A[0]), .Y(n4) );
  AND2X4 U4 ( .A(A[8]), .B(carry[8]), .Y(n2) );
  CLKAND2X8 U5 ( .A(A[6]), .B(carry[6]), .Y(n3) );
  INVXL U6 ( .A(n4), .Y(SUM[0]) );
  XOR2XL U7 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XOR2X4 U8 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  XOR2XL U9 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U10 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  CLKINVX8 U11 ( .A(n5), .Y(carry[3]) );
endmodule


module PWMConvert_DW01_inc_3 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [16:3] carry;

  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_14 ( .A(A[14]), .B(n3), .CO(carry[15]), .S(SUM[14]) );
  ADDHX4 U1_1_2 ( .A(A[2]), .B(n4), .CO(carry[3]), .S(SUM[2]) );
  ADDHX2 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(n2), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX4 U1_1_4 ( .A(A[4]), .B(n5), .CO(carry[5]), .S(SUM[4]) );
  CLKAND2X8 U1 ( .A(A[3]), .B(carry[3]), .Y(n5) );
  INVX6 U2 ( .A(n6), .Y(carry[11]) );
  BUFX6 U3 ( .A(A[0]), .Y(n1) );
  AND2X8 U4 ( .A(A[8]), .B(carry[8]), .Y(n2) );
  NAND2X4 U5 ( .A(A[10]), .B(carry[10]), .Y(n6) );
  NAND2X1 U6 ( .A(n8), .B(n9), .Y(SUM[13]) );
  NAND2X1 U7 ( .A(A[13]), .B(n16), .Y(n8) );
  NAND2X1 U8 ( .A(n7), .B(carry[13]), .Y(n9) );
  NAND2X1 U9 ( .A(carry[16]), .B(n13), .Y(n14) );
  AND2X2 U10 ( .A(carry[12]), .B(n12), .Y(n3) );
  AND2X2 U11 ( .A(A[1]), .B(n1), .Y(n4) );
  CLKINVX1 U12 ( .A(n16), .Y(carry[13]) );
  NAND2X1 U13 ( .A(A[12]), .B(carry[12]), .Y(n16) );
  CLKINVX1 U14 ( .A(n11), .Y(carry[16]) );
  NAND2X2 U15 ( .A(A[15]), .B(carry[15]), .Y(n11) );
  XOR2XL U16 ( .A(A[10]), .B(carry[10]), .Y(SUM[10]) );
  CLKINVX1 U17 ( .A(A[13]), .Y(n7) );
  XOR2XL U18 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  INVX8 U19 ( .A(n10), .Y(carry[7]) );
  NAND2X8 U20 ( .A(A[6]), .B(carry[6]), .Y(n10) );
  XOR2XL U21 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  AND2X2 U22 ( .A(A[12]), .B(A[13]), .Y(n12) );
  XOR2XL U23 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U24 ( .A(A[1]), .B(n1), .Y(SUM[1]) );
  XOR2XL U25 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  NAND2X1 U26 ( .A(n11), .B(A[16]), .Y(n15) );
  NAND2X1 U27 ( .A(n14), .B(n15), .Y(SUM[16]) );
  CLKINVX1 U28 ( .A(A[16]), .Y(n13) );
  XOR2XL U29 ( .A(A[3]), .B(carry[3]), .Y(SUM[3]) );
  CLKINVX1 U30 ( .A(n1), .Y(SUM[0]) );
endmodule


module PWMConvert_DW01_inc_4 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [16:2] carry;

  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(n4), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(n1), .B(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDHX2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHX4 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_15 ( .A(A[15]), .B(n3), .CO(carry[16]), .S(SUM[15]) );
  BUFX6 U1 ( .A(A[1]), .Y(n1) );
  INVX6 U2 ( .A(n5), .Y(carry[7]) );
  AND2X2 U3 ( .A(A[14]), .B(carry[14]), .Y(n3) );
  BUFX4 U4 ( .A(A[0]), .Y(n2) );
  AND2X4 U5 ( .A(A[2]), .B(carry[2]), .Y(n4) );
  XOR2X4 U6 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  INVXL U7 ( .A(n2), .Y(SUM[0]) );
  XOR2XL U8 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  NAND2X6 U9 ( .A(A[6]), .B(carry[6]), .Y(n5) );
  XOR2X1 U10 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2XL U11 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  CLKINVX8 U12 ( .A(n6), .Y(carry[9]) );
  NAND2X4 U13 ( .A(A[8]), .B(carry[8]), .Y(n6) );
  XOR2XL U14 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
endmodule


module PWMConvert_DW01_inc_5 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11;
  wire   [15:2] carry;

  ADDHX4 U1_1_14 ( .A(A[14]), .B(n2), .CO(carry[15]), .S(SUM[14]) );
  ADDHX4 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHX1 U1_1_4 ( .A(A[4]), .B(n3), .CO(carry[5]), .S(SUM[4]) );
  ADDHX2 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(n7), .CO(carry[8]), .S(SUM[7]) );
  CMPR22X2 U1_1_11 ( .A(A[11]), .B(n6), .CO(carry[12]), .S(SUM[11]) );
  NOR2X4 U1 ( .A(n10), .B(n8), .Y(n6) );
  XOR2X2 U2 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  XOR2X4 U3 ( .A(n4), .B(A[16]), .Y(SUM[16]) );
  BUFX8 U4 ( .A(A[0]), .Y(n1) );
  NAND2X6 U5 ( .A(A[8]), .B(carry[8]), .Y(n10) );
  AND2X2 U6 ( .A(A[12]), .B(carry[12]), .Y(n9) );
  CLKINVX4 U7 ( .A(n11), .Y(carry[2]) );
  NAND2X2 U8 ( .A(A[1]), .B(n1), .Y(n11) );
  AND2X2 U9 ( .A(A[6]), .B(carry[6]), .Y(n7) );
  NAND2X1 U10 ( .A(A[9]), .B(A[10]), .Y(n8) );
  AND2X2 U11 ( .A(A[13]), .B(n9), .Y(n2) );
  AND2X2 U12 ( .A(A[3]), .B(carry[3]), .Y(n3) );
  AND2X2 U13 ( .A(A[15]), .B(carry[15]), .Y(n4) );
  AND2X2 U14 ( .A(A[9]), .B(carry[9]), .Y(n5) );
  INVX1 U15 ( .A(n10), .Y(carry[9]) );
  XOR2XL U16 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XOR2XL U17 ( .A(A[10]), .B(n5), .Y(SUM[10]) );
  XOR2XL U18 ( .A(A[9]), .B(carry[9]), .Y(SUM[9]) );
  XOR2XL U19 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U20 ( .A(A[1]), .B(n1), .Y(SUM[1]) );
  XOR2XL U21 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XOR2X1 U22 ( .A(A[13]), .B(n9), .Y(SUM[13]) );
  XOR2XL U23 ( .A(A[3]), .B(carry[3]), .Y(SUM[3]) );
  CLKINVX1 U24 ( .A(n1), .Y(SUM[0]) );
endmodule


module PWMConvert_DW01_inc_6 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12;
  wire   [16:4] carry;

  ADDHX2 U1_1_14 ( .A(A[14]), .B(n2), .CO(carry[15]), .S(SUM[14]) );
  ADDHX1 U1_1_12 ( .A(A[12]), .B(n3), .CO(carry[13]), .S(SUM[12]) );
  ADDHX1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHX4 U1_1_3 ( .A(A[3]), .B(n6), .CO(carry[4]), .S(SUM[3]) );
  NAND2X8 U1 ( .A(A[6]), .B(n7), .Y(n12) );
  CLKAND2X12 U2 ( .A(A[5]), .B(carry[5]), .Y(n7) );
  CLKAND2X12 U3 ( .A(A[2]), .B(n4), .Y(n6) );
  XOR2X4 U4 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  AND2X2 U5 ( .A(A[1]), .B(A[0]), .Y(n4) );
  AND2X2 U6 ( .A(A[10]), .B(n1), .Y(n10) );
  XOR2X1 U7 ( .A(A[11]), .B(n11), .Y(SUM[11]) );
  AND2X2 U8 ( .A(A[9]), .B(n9), .Y(n1) );
  AND2X2 U9 ( .A(A[13]), .B(carry[13]), .Y(n2) );
  AND2X2 U10 ( .A(A[11]), .B(n10), .Y(n3) );
  NAND2X1 U11 ( .A(A[7]), .B(A[8]), .Y(n5) );
  NOR2X2 U12 ( .A(n12), .B(n5), .Y(n9) );
  AND2X2 U13 ( .A(A[7]), .B(carry[7]), .Y(n8) );
  INVX1 U14 ( .A(n12), .Y(carry[7]) );
  AND2XL U15 ( .A(A[10]), .B(n1), .Y(n11) );
  XOR2XL U16 ( .A(A[8]), .B(n8), .Y(SUM[8]) );
  XOR2XL U17 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  XOR2XL U18 ( .A(A[6]), .B(n7), .Y(SUM[6]) );
  XOR2XL U19 ( .A(A[9]), .B(n9), .Y(SUM[9]) );
  XOR2XL U20 ( .A(A[1]), .B(A[0]), .Y(SUM[1]) );
  XOR2XL U21 ( .A(A[10]), .B(n1), .Y(SUM[10]) );
  XOR2XL U22 ( .A(A[2]), .B(n4), .Y(SUM[2]) );
  XOR2XL U23 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  XOR2XL U24 ( .A(A[13]), .B(carry[13]), .Y(SUM[13]) );
  CLKINVX1 U25 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module PWMConvert_DW01_inc_7 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [16:2] carry;

  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(n3), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_13 ( .A(A[13]), .B(n4), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  CMPR22X4 U1_1_7 ( .A(A[7]), .B(n5), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(A[1]), .B(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDHX4 U1_1_9 ( .A(A[9]), .B(n2), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  CMPR22X2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  BUFX8 U1 ( .A(A[0]), .Y(n1) );
  INVXL U2 ( .A(n1), .Y(SUM[0]) );
  AND2X2 U3 ( .A(A[8]), .B(carry[8]), .Y(n2) );
  AND2X2 U4 ( .A(A[2]), .B(carry[2]), .Y(n3) );
  AND2X2 U5 ( .A(A[12]), .B(carry[12]), .Y(n4) );
  AND2X2 U6 ( .A(A[6]), .B(carry[6]), .Y(n5) );
  XOR2XL U7 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XOR2XL U8 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XOR2XL U9 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X4 U10 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  XOR2XL U11 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
endmodule


module PWMConvert_DW01_inc_8 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [16:2] carry;

  ADDHX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(n1), .B(n3), .CO(carry[2]), .S(SUM[1]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(n2), .CO(carry[16]), .S(SUM[15]) );
  CMPR22X2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  CMPR22X2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  BUFX8 U1 ( .A(A[1]), .Y(n1) );
  BUFX4 U2 ( .A(A[0]), .Y(n3) );
  AND2X4 U3 ( .A(A[14]), .B(carry[14]), .Y(n2) );
  XOR2X4 U4 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  INVXL U5 ( .A(n3), .Y(SUM[0]) );
  XOR2XL U6 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  INVX8 U7 ( .A(n4), .Y(carry[7]) );
  NAND2X6 U8 ( .A(A[6]), .B(carry[6]), .Y(n4) );
  XOR2X1 U9 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2XL U10 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  CLKINVX8 U11 ( .A(n5), .Y(carry[9]) );
  NAND2X4 U12 ( .A(A[8]), .B(carry[8]), .Y(n5) );
  XOR2XL U13 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  CLKINVX8 U14 ( .A(n6), .Y(carry[3]) );
  NAND2X6 U15 ( .A(A[2]), .B(carry[2]), .Y(n6) );
endmodule


module PWMConvert_DW01_inc_9 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
;
  wire   [15:4] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHX4 U1_1_14 ( .A(A[14]), .B(n10), .CO(carry[15]), .S(SUM[14]) );
  CMPR22X4 U1_1_12 ( .A(A[12]), .B(n7), .CO(carry[13]), .S(SUM[12]) );
  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_3 ( .A(A[3]), .B(n15), .CO(carry[4]), .S(SUM[3]) );
  CLKAND2X8 U1 ( .A(A[2]), .B(n3), .Y(n15) );
  BUFX8 U2 ( .A(A[0]), .Y(n1) );
  INVXL U3 ( .A(n1), .Y(SUM[0]) );
  CLKAND2X6 U4 ( .A(A[1]), .B(n1), .Y(n3) );
  CLKAND2X12 U5 ( .A(A[11]), .B(n8), .Y(n7) );
  AND2X2 U6 ( .A(A[13]), .B(carry[13]), .Y(n10) );
  AND2X2 U7 ( .A(A[9]), .B(n11), .Y(n13) );
  AND2X2 U8 ( .A(n5), .B(n6), .Y(n11) );
  AND2X2 U9 ( .A(carry[6]), .B(A[6]), .Y(n5) );
  AND2X2 U10 ( .A(A[6]), .B(carry[6]), .Y(n16) );
  AND2X2 U11 ( .A(A[10]), .B(n13), .Y(n8) );
  XOR2X1 U12 ( .A(n2), .B(A[16]), .Y(SUM[16]) );
  AND2X2 U13 ( .A(A[15]), .B(carry[15]), .Y(n2) );
  AND2X2 U14 ( .A(A[7]), .B(n16), .Y(n4) );
  XOR2XL U15 ( .A(A[1]), .B(n1), .Y(SUM[1]) );
  AND2X2 U16 ( .A(A[8]), .B(A[7]), .Y(n6) );
  AND2XL U17 ( .A(A[10]), .B(n13), .Y(n9) );
  XOR2X4 U18 ( .A(A[15]), .B(carry[15]), .Y(SUM[15]) );
  XOR2XL U19 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  XOR2X1 U20 ( .A(A[10]), .B(n14), .Y(SUM[10]) );
  AND2XL U21 ( .A(A[8]), .B(n4), .Y(n12) );
  XOR2XL U22 ( .A(A[8]), .B(n4), .Y(SUM[8]) );
  XOR2X1 U23 ( .A(A[9]), .B(n12), .Y(SUM[9]) );
  AND2XL U24 ( .A(A[9]), .B(n12), .Y(n14) );
  XOR2XL U25 ( .A(A[11]), .B(n9), .Y(SUM[11]) );
  XOR2XL U26 ( .A(A[2]), .B(n3), .Y(SUM[2]) );
  XOR2XL U27 ( .A(A[13]), .B(carry[13]), .Y(SUM[13]) );
endmodule


module PWMConvert_DW01_inc_10 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [13:3] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(n9), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(n8), .CO(carry[5]), .S(SUM[4]) );
  ADDHX4 U1_1_12 ( .A(A[12]), .B(n2), .CO(carry[13]), .S(SUM[12]) );
  BUFX8 U1 ( .A(A[0]), .Y(n1) );
  INVXL U2 ( .A(n1), .Y(SUM[0]) );
  CLKAND2X8 U3 ( .A(A[1]), .B(n1), .Y(n7) );
  NAND2X2 U4 ( .A(n12), .B(n13), .Y(SUM[14]) );
  NOR2X2 U5 ( .A(n24), .B(n14), .Y(n18) );
  NAND2X1 U6 ( .A(A[3]), .B(A[4]), .Y(n14) );
  NAND2X1 U7 ( .A(A[2]), .B(n7), .Y(n24) );
  CLKINVX1 U8 ( .A(n5), .Y(n11) );
  CLKINVX1 U9 ( .A(n24), .Y(carry[3]) );
  AND2X2 U10 ( .A(A[7]), .B(n21), .Y(n16) );
  NAND2X1 U11 ( .A(n10), .B(n5), .Y(n13) );
  NAND2X1 U12 ( .A(A[14]), .B(n11), .Y(n12) );
  XOR2X1 U13 ( .A(n3), .B(A[16]), .Y(SUM[16]) );
  AND2X2 U14 ( .A(A[11]), .B(n4), .Y(n2) );
  AND2X2 U15 ( .A(A[15]), .B(n6), .Y(n3) );
  AND2X2 U16 ( .A(A[10]), .B(n22), .Y(n4) );
  AND2X2 U17 ( .A(A[13]), .B(carry[13]), .Y(n5) );
  AND2X2 U18 ( .A(carry[13]), .B(n15), .Y(n6) );
  AND2X2 U19 ( .A(A[3]), .B(carry[3]), .Y(n8) );
  CLKAND2X12 U20 ( .A(A[5]), .B(n18), .Y(n9) );
  CLKINVX1 U21 ( .A(A[14]), .Y(n10) );
  XOR2X2 U22 ( .A(A[15]), .B(n6), .Y(SUM[15]) );
  AND2X2 U23 ( .A(A[13]), .B(A[14]), .Y(n15) );
  AND2X2 U24 ( .A(A[8]), .B(n16), .Y(n19) );
  AND2X1 U25 ( .A(A[9]), .B(n20), .Y(n23) );
  AND2X2 U26 ( .A(A[6]), .B(n9), .Y(n21) );
  AND2XL U27 ( .A(A[7]), .B(n21), .Y(n17) );
  XOR2XL U28 ( .A(A[5]), .B(carry[5]), .Y(SUM[5]) );
  AND2X2 U29 ( .A(A[9]), .B(n19), .Y(n22) );
  AND2XL U30 ( .A(A[8]), .B(n17), .Y(n20) );
  XOR2XL U31 ( .A(A[3]), .B(carry[3]), .Y(SUM[3]) );
  XOR2XL U32 ( .A(A[1]), .B(n1), .Y(SUM[1]) );
  XOR2XL U33 ( .A(A[8]), .B(n17), .Y(SUM[8]) );
  XOR2XL U34 ( .A(A[11]), .B(n4), .Y(SUM[11]) );
  XOR2X1 U35 ( .A(A[10]), .B(n23), .Y(SUM[10]) );
  XOR2XL U36 ( .A(A[7]), .B(carry[7]), .Y(SUM[7]) );
  XOR2XL U37 ( .A(A[9]), .B(n20), .Y(SUM[9]) );
  XOR2XL U38 ( .A(A[2]), .B(n7), .Y(SUM[2]) );
  XOR2XL U39 ( .A(A[13]), .B(carry[13]), .Y(SUM[13]) );
endmodule


module PWMConvert_DW01_inc_11 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [16:2] carry;

  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(n4), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(n1), .B(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDHX2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHX4 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_15 ( .A(A[15]), .B(n3), .CO(carry[16]), .S(SUM[15]) );
  BUFX6 U1 ( .A(A[1]), .Y(n1) );
  INVX6 U2 ( .A(n5), .Y(carry[7]) );
  AND2X2 U3 ( .A(A[14]), .B(carry[14]), .Y(n3) );
  BUFX4 U4 ( .A(A[0]), .Y(n2) );
  AND2X4 U5 ( .A(A[2]), .B(carry[2]), .Y(n4) );
  XOR2X4 U6 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  INVXL U7 ( .A(n2), .Y(SUM[0]) );
  XOR2XL U8 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  NAND2X6 U9 ( .A(A[6]), .B(carry[6]), .Y(n5) );
  XOR2X1 U10 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2XL U11 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  CLKINVX8 U12 ( .A(n6), .Y(carry[9]) );
  NAND2X4 U13 ( .A(A[8]), .B(carry[8]), .Y(n6) );
  XOR2XL U14 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
endmodule


module PWMConvert_DW01_inc_12 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [16:2] carry;

  ADDHX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(n1), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(n2), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  CMPR22X2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  CMPR22X2 U1_1_1 ( .A(A[1]), .B(n3), .CO(carry[2]), .S(SUM[1]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHX2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  BUFX4 U1 ( .A(A[0]), .Y(n3) );
  AND2X4 U2 ( .A(A[8]), .B(carry[8]), .Y(n1) );
  CLKAND2X8 U3 ( .A(A[6]), .B(carry[6]), .Y(n2) );
  INVXL U4 ( .A(n3), .Y(SUM[0]) );
  XOR2XL U5 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XOR2X4 U6 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  XOR2XL U7 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2XL U8 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  CLKINVX8 U9 ( .A(n4), .Y(carry[3]) );
  NAND2X6 U10 ( .A(A[2]), .B(carry[2]), .Y(n4) );
endmodule


module PWMConvert_DW01_inc_13 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [16:2] carry;

  ADDHX1 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(n1), .B(n3), .CO(carry[2]), .S(SUM[1]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(n2), .CO(carry[16]), .S(SUM[15]) );
  CMPR22X2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  CMPR22X2 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  XOR2X2 U1 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  BUFX8 U2 ( .A(A[1]), .Y(n1) );
  BUFX4 U3 ( .A(A[0]), .Y(n3) );
  AND2X4 U4 ( .A(A[14]), .B(carry[14]), .Y(n2) );
  INVXL U5 ( .A(n3), .Y(SUM[0]) );
  XOR2XL U6 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  INVX8 U7 ( .A(n4), .Y(carry[7]) );
  NAND2X6 U8 ( .A(A[6]), .B(carry[6]), .Y(n4) );
  XOR2X1 U9 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2XL U10 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  CLKINVX8 U11 ( .A(n5), .Y(carry[9]) );
  NAND2X4 U12 ( .A(A[8]), .B(carry[8]), .Y(n5) );
  XOR2XL U13 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
  CLKINVX8 U14 ( .A(n6), .Y(carry[3]) );
  NAND2X6 U15 ( .A(A[2]), .B(carry[2]), .Y(n6) );
endmodule


module PWMConvert_DW01_inc_14 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5, n6;
  wire   [16:2] carry;

  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(n4), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(n1), .B(n2), .CO(carry[2]), .S(SUM[1]) );
  ADDHX2 U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHX4 U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHX1 U1_1_15 ( .A(A[15]), .B(n3), .CO(carry[16]), .S(SUM[15]) );
  BUFX6 U1 ( .A(A[1]), .Y(n1) );
  INVX6 U2 ( .A(n5), .Y(carry[7]) );
  AND2X2 U3 ( .A(A[14]), .B(carry[14]), .Y(n3) );
  BUFX4 U4 ( .A(A[0]), .Y(n2) );
  AND2X4 U5 ( .A(A[2]), .B(carry[2]), .Y(n4) );
  XOR2X4 U6 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  INVXL U7 ( .A(n2), .Y(SUM[0]) );
  XOR2XL U8 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  NAND2X6 U9 ( .A(A[6]), .B(carry[6]), .Y(n5) );
  XOR2X1 U10 ( .A(A[14]), .B(carry[14]), .Y(SUM[14]) );
  XOR2XL U11 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  CLKINVX8 U12 ( .A(n6), .Y(carry[9]) );
  NAND2X4 U13 ( .A(A[8]), .B(carry[8]), .Y(n6) );
  XOR2XL U14 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
endmodule


module PWMConvert_DW01_inc_15 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n4, n5;
  wire   [16:2] carry;

  ADDHX2 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  CMPR22X4 U1_1_3 ( .A(A[3]), .B(n3), .CO(carry[4]), .S(SUM[3]) );
  CMPR22X4 U1_1_13 ( .A(A[13]), .B(n4), .CO(carry[14]), .S(SUM[13]) );
  ADDHX4 U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  CMPR22X4 U1_1_7 ( .A(A[7]), .B(n5), .CO(carry[8]), .S(SUM[7]) );
  ADDHX4 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHX4 U1_1_1 ( .A(A[1]), .B(n1), .CO(carry[2]), .S(SUM[1]) );
  ADDHX4 U1_1_9 ( .A(A[9]), .B(n2), .CO(carry[10]), .S(SUM[9]) );
  ADDHX4 U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  CMPR22X2 U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHX4 U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  BUFX8 U1 ( .A(A[0]), .Y(n1) );
  INVXL U2 ( .A(n1), .Y(SUM[0]) );
  AND2X2 U3 ( .A(A[8]), .B(carry[8]), .Y(n2) );
  AND2X2 U4 ( .A(A[2]), .B(carry[2]), .Y(n3) );
  AND2X2 U5 ( .A(A[12]), .B(carry[12]), .Y(n4) );
  AND2X2 U6 ( .A(A[6]), .B(carry[6]), .Y(n5) );
  XOR2XL U7 ( .A(A[6]), .B(carry[6]), .Y(SUM[6]) );
  XOR2XL U8 ( .A(A[12]), .B(carry[12]), .Y(SUM[12]) );
  XOR2XL U9 ( .A(A[8]), .B(carry[8]), .Y(SUM[8]) );
  XOR2X4 U10 ( .A(carry[16]), .B(A[16]), .Y(SUM[16]) );
  XOR2XL U11 ( .A(A[2]), .B(carry[2]), .Y(SUM[2]) );
endmodule


module PWMConvert_DW01_inc_16 ( A, SUM );
  input [10:0] A;
  output [10:0] SUM;
  wire   n1, n2, n3, n4;
  wire   [10:2] carry;

  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHX1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  ADDHX2 U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHX1 U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHX1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHX1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  NAND2X2 U1 ( .A(n3), .B(n4), .Y(SUM[10]) );
  NAND2X2 U2 ( .A(n1), .B(A[10]), .Y(n4) );
  NAND2X1 U3 ( .A(carry[10]), .B(n2), .Y(n3) );
  INVX2 U4 ( .A(carry[10]), .Y(n1) );
  CLKINVX1 U5 ( .A(A[10]), .Y(n2) );
  CLKINVX1 U6 ( .A(A[0]), .Y(SUM[0]) );
endmodule


module PWMConvert ( GCK, Vsync, mode, rst, OUT, data, addr, en );
  output [15:0] OUT;
  input [15:0] data;
  output [8:0] addr;
  input GCK, Vsync, mode, rst;
  output en;
  wire   r_push_reg, N39, N40, N41, N42, N43, N45, N48, N49, N50, N51, N52,
         N53, N54, N55, N56, N57, N58, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126,
         N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137,
         N138, N139, N140, N141, N142, N143, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N210, N211, N212, N213,
         N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393,
         N410, N411, N412, N413, N414, N415, N416, N417, N418, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N428, N429, N430, N431,
         N432, N433, N434, N435, N436, N437, N438, N439, N440, N441, N442,
         N443, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N510, N511, N512, N513, N514, N515, N516, N517, N518,
         N519, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N536, N537, N538, N539, N540,
         N541, N542, N543, N560, N561, N562, N563, N564, N565, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589,
         N590, N591, N592, N593, N610, N611, N612, N613, N614, N615, N616,
         N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627,
         N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638,
         N639, N640, N641, N642, N643, N660, N661, N662, N663, N664, N665,
         N666, N667, N668, N669, N670, N671, N672, N673, N674, N675, N676,
         N677, N678, N679, N680, N681, N682, N683, N684, N685, N686, N687,
         N688, N689, N690, N691, N692, N693, N710, N711, N712, N713, N714,
         N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725,
         N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N760, N761, N762, N763,
         N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N810, N811, N812,
         N813, N814, N815, N816, N817, N818, N819, N820, N821, N822, N823,
         N824, N825, N826, N827, N828, N829, N830, N831, N832, N833, N834,
         N835, N836, N837, N838, N839, N840, N841, N842, N843, N860, N861,
         N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872,
         N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883,
         N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n47, n63, n79, n95, n1110, n2740,
         n2750, n2800, n2810, n8120, n8130, n8140, n8150, n8160, n8170, n8180,
         n8190, n8200, n8210, n8220, n8230, n8240, n8250, n8260, n8280, n8290,
         n8300, n8310, n8320, n8330, n8340, n8350, n8360, n8370, n8380, n8390,
         n8400, n8410, n8420, n8430, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n8600, n8610,
         n8620, n8630, n8640, n8650, n8660, n8670, n8680, n8690, n8700, n8710,
         n8720, n8730, n8740, n8750, n8760, n8770, n8780, n8790, n8800, n8810,
         n8820, n8830, n8840, n8850, n8860, n8870, n8880, n8890, n8900, n8910,
         n8920, n8930, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1075, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         N9070, N9060, N9050, N9040, N9030, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n1830, n1840, n1900, n1910, n1920, n1930,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n3600, n3610, n3620, n3630, n3640, n3650,
         n3660, n3670, n3680, n3690, n3700, n3710, n3720, n3730, n3740, n3750,
         n3760, n3770, n3780, n3790, n3800, n3810, n3820, n3830, n3840, n3850,
         n3860, n3870, n3880, n3890, n3900, n3910, n3920, n3930, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n4100, n4110, n4120, n4130, n4140, n4150, n4160,
         n4170, n4180, n4190, n4200, n4210, n4220, n4230, n4240, n4250, n4260,
         n4270, n4280, n4290, n4300, n4310, n4320, n4330, n4340, n4350, n4360,
         n4370, n4380, n4390, n4400, n4410, n4420, n4430, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n4600, n4610, n4620, n4630, n4640, n4650, n4660, n4670,
         n4680, n4690, n4700, n4710, n4720, n4730, n4740, n4750, n4760, n4770,
         n4780, n4790, n4800, n4810, n4820, n4830, n4840, n4850, n4860, n4870,
         n4880, n4890, n4900, n4910, n4920, n4930, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n5100, n5110, n5120, n5130, n5140, n5150, n5160, n5170, n5180,
         n5190, n5200, n5210, n5220, n5230, n5240, n5250, n5260, n5270, n5280,
         n5290, n5300, n5310, n5320, n5330, n5340, n5350, n5360, n5370, n5380,
         n5390, n5400, n5410, n5420, n5430, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n5600,
         n5610, n5620, n5630, n5640, n5650, n5660, n5670, n5680, n5690, n5700,
         n5710, n5720, n5730, n5740, n5750, n5760, n5770, n5780, n5790, n5800,
         n5810, n5820, n5830, n5840, n5850, n5860, n5870, n5880, n5890, n5900,
         n5910, n5920, n5930, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n6100, n6110, n6120,
         n6130, n6140, n6150, n6160, n6170, n6180, n6190, n6200, n6210, n6220,
         n6230, n6240, n6250, n6260, n6270, n6280, n6290, n6300, n6310, n6320,
         n6330, n6340, n6350, n6360, n6370, n6380, n6390, n6400, n6410, n6420,
         n6430, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n6600, n6610, n6620, n6630, n6640,
         n6650, n6660, n6670, n6680, n6690, n6700, n6710, n6720, n6730, n6740,
         n6750, n6760, n6770, n6780, n6790, n6800, n6810, n6820, n6830, n6840,
         n6850, n6860, n6870, n6880, n6890, n6900, n6910, n6920, n6930, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n7100, n7110, n7120, n7130, n7140, n7150,
         n7160, n7170, n7180, n7190, n7200, n7210, n7220, n7230, n7240, n7250,
         n7260, n7270, n7280, n7290, n7300, n7310, n7320, n7330, n7340, n7350,
         n7360, n7370, n7380, n7390, n7400, n7410, n7420, n7430, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n7600, n7610, n7620, n7630, n7640, n7650, n7660,
         n7670, n7680, n7690, n7700, n7710, n7720, n7730, n7740, n7750, n7760,
         n7770, n7780, n7790, n7800, n7810, n7820, n7830, n7840, n7850, n7860,
         n7870, n7880, n7890, n7900, n7910, n7920, n7930, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n8100, n8110, n8270, n1019;
  wire   [2:0] out_cs;
  wire   [4:0] cnt;
  wire   [10:9] rd_addr;
  wire   [254:0] rd_reg;
  wire   [255:0] out_buffer;
  wire   [4:2] add_101_aco_carry;

  DFFRX1 rd_reg_reg_15__5_ ( .D(n907), .CK(GCK), .RN(n4390), .Q(rd_reg[5]), 
        .QN(n87) );
  DFFRX1 rd_reg_reg_15__4_ ( .D(n8910), .CK(GCK), .RN(n4370), .Q(rd_reg[4]), 
        .QN(n94) );
  DFFRX1 rd_reg_reg_15__3_ ( .D(n8750), .CK(GCK), .RN(n4370), .Q(rd_reg[3]), 
        .QN(n91) );
  DFFRX1 rd_reg_reg_15__2_ ( .D(n859), .CK(GCK), .RN(n4410), .Q(rd_reg[2]), 
        .QN(n93) );
  DFFRX1 rd_reg_reg_15__1_ ( .D(n8430), .CK(GCK), .RN(n4360), .Q(rd_reg[1]), 
        .QN(n92) );
  DFFRX1 rd_reg_reg_15__0_ ( .D(n5860), .CK(GCK), .RN(n4360), .Q(rd_reg[0]) );
  DFFRX1 rd_reg_reg_15__12_ ( .D(n5830), .CK(GCK), .RN(n4420), .Q(rd_reg[12]), 
        .QN(n103) );
  DFFRX1 rd_reg_reg_15__11_ ( .D(n1003), .CK(GCK), .RN(n4410), .Q(rd_reg[11]), 
        .QN(n102) );
  DFFRX1 rd_reg_reg_15__10_ ( .D(n987), .CK(GCK), .RN(n4400), .Q(rd_reg[10]), 
        .QN(n101) );
  DFFRX1 rd_reg_reg_15__9_ ( .D(n971), .CK(GCK), .RN(n4400), .Q(rd_reg[9]), 
        .QN(n100) );
  DFFRX1 rd_reg_reg_15__8_ ( .D(n955), .CK(GCK), .RN(n4390), .Q(rd_reg[8]), 
        .QN(n99) );
  DFFRX1 rd_reg_reg_15__7_ ( .D(n939), .CK(GCK), .RN(n4380), .Q(rd_reg[7]), 
        .QN(n98) );
  DFFRX1 rd_reg_reg_15__6_ ( .D(n923), .CK(GCK), .RN(n4380), .Q(rd_reg[6]), 
        .QN(n104) );
  DFFRX1 rd_reg_reg_15__13_ ( .D(n5840), .CK(GCK), .RN(n4420), .Q(rd_reg[13]), 
        .QN(n97) );
  DFFRX1 rd_reg_reg_15__14_ ( .D(n1051), .CK(GCK), .RN(n4350), .Q(rd_reg[14]), 
        .QN(n105) );
  DFFRX1 r_carry_60_reg ( .D(n1080), .CK(GCK), .RN(n400), .Q(n5180) );
  DFFRX1 out_buffer_reg_15__10_ ( .D(N887), .CK(GCK), .RN(n402), .Q(
        out_buffer[10]) );
  DFFRX1 out_buffer_reg_15__11_ ( .D(N888), .CK(GCK), .RN(n402), .Q(
        out_buffer[11]) );
  DFFRX1 out_buffer_reg_15__13_ ( .D(N890), .CK(GCK), .RN(n402), .Q(
        out_buffer[13]) );
  DFFRX1 out_buffer_reg_15__14_ ( .D(N891), .CK(GCK), .RN(n402), .Q(
        out_buffer[14]) );
  DFFRX1 out_buffer_reg_15__15_ ( .D(N892), .CK(GCK), .RN(n402), .Q(
        out_buffer[15]) );
  DFFRX1 out_buffer_reg_13__10_ ( .D(N787), .CK(GCK), .RN(n404), .Q(
        out_buffer[42]) );
  DFFRX1 out_buffer_reg_13__11_ ( .D(N788), .CK(GCK), .RN(n405), .Q(
        out_buffer[43]) );
  DFFRX1 out_buffer_reg_13__12_ ( .D(N789), .CK(GCK), .RN(n405), .Q(
        out_buffer[44]) );
  DFFRX1 out_buffer_reg_13__13_ ( .D(N790), .CK(GCK), .RN(n405), .Q(
        out_buffer[45]) );
  DFFRX1 out_buffer_reg_13__14_ ( .D(N791), .CK(GCK), .RN(n405), .Q(
        out_buffer[46]) );
  DFFRX1 out_buffer_reg_13__15_ ( .D(N792), .CK(GCK), .RN(n405), .Q(
        out_buffer[47]) );
  DFFRX1 out_buffer_reg_12__11_ ( .D(N738), .CK(GCK), .RN(n406), .Q(
        out_buffer[59]) );
  DFFRX1 out_buffer_reg_12__14_ ( .D(N741), .CK(GCK), .RN(n406), .Q(
        out_buffer[62]) );
  DFFRX1 out_buffer_reg_11__10_ ( .D(N687), .CK(GCK), .RN(n407), .Q(
        out_buffer[74]) );
  DFFRX1 out_buffer_reg_11__11_ ( .D(N688), .CK(GCK), .RN(n407), .Q(
        out_buffer[75]) );
  DFFRX1 out_buffer_reg_11__12_ ( .D(N689), .CK(GCK), .RN(n407), .Q(
        out_buffer[76]) );
  DFFRX1 out_buffer_reg_11__13_ ( .D(N690), .CK(GCK), .RN(n408), .Q(
        out_buffer[77]) );
  DFFRX1 out_buffer_reg_11__15_ ( .D(N692), .CK(GCK), .RN(n408), .Q(
        out_buffer[79]) );
  DFFRX1 out_buffer_reg_10__11_ ( .D(N638), .CK(GCK), .RN(n409), .Q(
        out_buffer[91]) );
  DFFRX1 out_buffer_reg_10__14_ ( .D(N641), .CK(GCK), .RN(n409), .Q(
        out_buffer[94]) );
  DFFRX1 out_buffer_reg_9__12_ ( .D(N589), .CK(GCK), .RN(n4100), .Q(
        out_buffer[108]) );
  DFFRX1 out_buffer_reg_9__14_ ( .D(N591), .CK(GCK), .RN(n4100), .Q(
        out_buffer[110]) );
  DFFRX1 out_buffer_reg_9__15_ ( .D(N592), .CK(GCK), .RN(n4110), .Q(
        out_buffer[111]) );
  DFFRX1 out_buffer_reg_8__10_ ( .D(N537), .CK(GCK), .RN(n4120), .Q(
        out_buffer[122]) );
  DFFRX1 out_buffer_reg_8__11_ ( .D(N538), .CK(GCK), .RN(n4120), .Q(
        out_buffer[123]) );
  DFFRX1 out_buffer_reg_8__13_ ( .D(N540), .CK(GCK), .RN(n4120), .Q(
        out_buffer[125]) );
  DFFRX1 out_buffer_reg_8__14_ ( .D(N541), .CK(GCK), .RN(n4120), .Q(
        out_buffer[126]) );
  DFFRX1 out_buffer_reg_7__10_ ( .D(N487), .CK(GCK), .RN(n4130), .Q(
        out_buffer[138]) );
  DFFRX1 out_buffer_reg_7__11_ ( .D(N488), .CK(GCK), .RN(n4130), .Q(
        out_buffer[139]) );
  DFFRX1 out_buffer_reg_7__12_ ( .D(N489), .CK(GCK), .RN(n4130), .Q(
        out_buffer[140]) );
  DFFRX1 out_buffer_reg_7__13_ ( .D(N490), .CK(GCK), .RN(n4130), .Q(
        out_buffer[141]) );
  DFFRX1 out_buffer_reg_7__15_ ( .D(N492), .CK(GCK), .RN(n4130), .Q(
        out_buffer[143]) );
  DFFRX1 out_buffer_reg_6__12_ ( .D(N439), .CK(GCK), .RN(n4150), .Q(
        out_buffer[156]) );
  DFFRX1 out_buffer_reg_6__14_ ( .D(N441), .CK(GCK), .RN(n4150), .Q(
        out_buffer[158]) );
  DFFRX1 out_buffer_reg_5__12_ ( .D(N389), .CK(GCK), .RN(n4160), .Q(
        out_buffer[172]) );
  DFFRX1 out_buffer_reg_4__11_ ( .D(N338), .CK(GCK), .RN(n4170), .Q(
        out_buffer[187]) );
  DFFRX1 out_buffer_reg_4__12_ ( .D(N339), .CK(GCK), .RN(n4170), .Q(
        out_buffer[188]) );
  DFFRX1 out_buffer_reg_4__13_ ( .D(N340), .CK(GCK), .RN(n4170), .Q(
        out_buffer[189]) );
  DFFRX1 out_buffer_reg_4__15_ ( .D(N342), .CK(GCK), .RN(n4180), .Q(
        out_buffer[191]) );
  DFFRX1 out_buffer_reg_3__10_ ( .D(N287), .CK(GCK), .RN(n4190), .Q(
        out_buffer[202]) );
  DFFRX1 out_buffer_reg_3__11_ ( .D(N288), .CK(GCK), .RN(n4190), .Q(
        out_buffer[203]) );
  DFFRX1 out_buffer_reg_3__12_ ( .D(N289), .CK(GCK), .RN(n4190), .Q(
        out_buffer[204]) );
  DFFRX1 out_buffer_reg_3__13_ ( .D(N290), .CK(GCK), .RN(n4190), .Q(
        out_buffer[205]) );
  DFFRX1 out_buffer_reg_3__14_ ( .D(N291), .CK(GCK), .RN(n4190), .Q(
        out_buffer[206]) );
  DFFRX1 out_buffer_reg_3__15_ ( .D(N292), .CK(GCK), .RN(n4190), .Q(
        out_buffer[207]) );
  DFFRX1 out_buffer_reg_2__10_ ( .D(N237), .CK(GCK), .RN(n4200), .Q(
        out_buffer[218]) );
  DFFRX1 out_buffer_reg_2__11_ ( .D(N238), .CK(GCK), .RN(n4200), .Q(
        out_buffer[219]) );
  DFFRX1 out_buffer_reg_2__12_ ( .D(N239), .CK(GCK), .RN(n4200), .Q(
        out_buffer[220]) );
  DFFRX1 out_buffer_reg_2__13_ ( .D(N240), .CK(GCK), .RN(n4200), .Q(
        out_buffer[221]) );
  DFFRX1 out_buffer_reg_2__15_ ( .D(N242), .CK(GCK), .RN(n4200), .Q(
        out_buffer[223]) );
  DFFRX1 out_buffer_reg_1__10_ ( .D(N187), .CK(GCK), .RN(n4210), .Q(
        out_buffer[234]) );
  DFFRX1 out_buffer_reg_1__11_ ( .D(N188), .CK(GCK), .RN(n4220), .Q(
        out_buffer[235]) );
  DFFRX1 out_buffer_reg_1__12_ ( .D(N189), .CK(GCK), .RN(n4220), .Q(
        out_buffer[236]) );
  DFFRX1 out_buffer_reg_1__13_ ( .D(N190), .CK(GCK), .RN(n4220), .Q(
        out_buffer[237]) );
  DFFRX1 out_buffer_reg_1__15_ ( .D(N192), .CK(GCK), .RN(n4220), .Q(
        out_buffer[239]) );
  DFFRX1 out_buffer_reg_0__10_ ( .D(N137), .CK(GCK), .RN(n4230), .Q(
        out_buffer[250]) );
  DFFRX1 out_buffer_reg_0__11_ ( .D(N138), .CK(GCK), .RN(n4230), .Q(
        out_buffer[251]) );
  DFFRX1 out_buffer_reg_0__13_ ( .D(N140), .CK(GCK), .RN(n4230), .Q(
        out_buffer[253]) );
  DFFRX1 out_buffer_reg_0__14_ ( .D(N141), .CK(GCK), .RN(n4230), .Q(
        out_buffer[254]) );
  DFFRX1 out_cs_reg_0_ ( .D(n1094), .CK(GCK), .RN(n399), .Q(out_cs[0]), .QN(
        n86) );
  DFFRX1 rd_addr_reg_9_ ( .D(n1082), .CK(GCK), .RN(n400), .Q(rd_addr[9]), .QN(
        n1080) );
  DFFRX1 rd_addr_reg_5_ ( .D(n1086), .CK(GCK), .RN(n400), .Q(addr[5]), .QN(n9)
         );
  DFFRX1 rd_addr_reg_6_ ( .D(n1085), .CK(GCK), .RN(n400), .Q(addr[6]), .QN(n10) );
  DFFRX1 rd_addr_reg_7_ ( .D(n1084), .CK(GCK), .RN(n400), .Q(addr[7]), .QN(n11) );
  DFFRX1 rd_addr_reg_8_ ( .D(n1083), .CK(GCK), .RN(n400), .Q(addr[8]), .QN(n12) );
  DFFSX1 rd_addr_reg_4_ ( .D(n1087), .CK(GCK), .SN(n4230), .Q(addr[4]), .QN(n8) );
  DFFRX2 OUT_reg_15_ ( .D(N893), .CK(GCK), .RN(n401), .Q(OUT[15]) );
  DFFRX2 OUT_reg_14_ ( .D(N843), .CK(GCK), .RN(n402), .Q(OUT[14]) );
  DFFRX2 OUT_reg_13_ ( .D(N793), .CK(GCK), .RN(n404), .Q(OUT[13]) );
  DFFRX2 OUT_reg_12_ ( .D(N743), .CK(GCK), .RN(n405), .Q(OUT[12]) );
  DFFRX2 OUT_reg_11_ ( .D(N693), .CK(GCK), .RN(n406), .Q(OUT[11]) );
  DFFRX2 OUT_reg_10_ ( .D(N643), .CK(GCK), .RN(n408), .Q(OUT[10]) );
  DFFRX2 OUT_reg_9_ ( .D(N593), .CK(GCK), .RN(n409), .Q(OUT[9]) );
  DFFRX2 OUT_reg_8_ ( .D(N543), .CK(GCK), .RN(n4110), .Q(OUT[8]) );
  DFFRX2 OUT_reg_7_ ( .D(N493), .CK(GCK), .RN(n4120), .Q(OUT[7]) );
  DFFRX2 OUT_reg_6_ ( .D(N443), .CK(GCK), .RN(n4130), .Q(OUT[6]) );
  DFFRX2 OUT_reg_5_ ( .D(N393), .CK(GCK), .RN(n4150), .Q(OUT[5]) );
  DFFRX2 OUT_reg_4_ ( .D(N343), .CK(GCK), .RN(n4160), .Q(OUT[4]) );
  DFFRX2 OUT_reg_3_ ( .D(N293), .CK(GCK), .RN(n4180), .Q(OUT[3]) );
  DFFRX2 OUT_reg_2_ ( .D(N243), .CK(GCK), .RN(n4190), .Q(OUT[2]) );
  DFFRX2 OUT_reg_1_ ( .D(N193), .CK(GCK), .RN(n4210), .Q(OUT[1]) );
  DFFRX2 OUT_reg_0_ ( .D(N143), .CK(GCK), .RN(n4220), .Q(OUT[0]) );
  DFFRX1 out_buffer_reg_15__5_ ( .D(N882), .CK(GCK), .RN(n401), .Q(
        out_buffer[5]) );
  DFFRX1 out_buffer_reg_15__7_ ( .D(N884), .CK(GCK), .RN(n401), .Q(
        out_buffer[7]) );
  DFFRX1 out_buffer_reg_15__9_ ( .D(N886), .CK(GCK), .RN(n402), .Q(
        out_buffer[9]) );
  DFFRX1 out_buffer_reg_14__7_ ( .D(N834), .CK(GCK), .RN(n403), .Q(
        out_buffer[23]) );
  DFFRX1 out_buffer_reg_13__4_ ( .D(N781), .CK(GCK), .RN(n404), .Q(
        out_buffer[36]) );
  DFFRX1 out_buffer_reg_13__5_ ( .D(N782), .CK(GCK), .RN(n404), .Q(
        out_buffer[37]) );
  DFFRX1 out_buffer_reg_13__7_ ( .D(N784), .CK(GCK), .RN(n404), .Q(
        out_buffer[39]) );
  DFFRX1 out_buffer_reg_13__9_ ( .D(N786), .CK(GCK), .RN(n404), .Q(
        out_buffer[41]) );
  DFFRX1 out_buffer_reg_12__4_ ( .D(N731), .CK(GCK), .RN(n405), .Q(
        out_buffer[52]) );
  DFFRX1 out_buffer_reg_12__5_ ( .D(N732), .CK(GCK), .RN(n405), .Q(
        out_buffer[53]) );
  DFFRX1 out_buffer_reg_12__7_ ( .D(N734), .CK(GCK), .RN(n406), .Q(
        out_buffer[55]) );
  DFFRX1 out_buffer_reg_12__9_ ( .D(N736), .CK(GCK), .RN(n406), .Q(
        out_buffer[57]) );
  DFFRX1 out_buffer_reg_11__4_ ( .D(N681), .CK(GCK), .RN(n407), .Q(
        out_buffer[68]) );
  DFFRX1 out_buffer_reg_11__5_ ( .D(N682), .CK(GCK), .RN(n407), .Q(
        out_buffer[69]) );
  DFFRX1 out_buffer_reg_11__7_ ( .D(N684), .CK(GCK), .RN(n407), .Q(
        out_buffer[71]) );
  DFFRX1 out_buffer_reg_11__9_ ( .D(N686), .CK(GCK), .RN(n407), .Q(
        out_buffer[73]) );
  DFFRX1 out_buffer_reg_10__4_ ( .D(N631), .CK(GCK), .RN(n408), .Q(
        out_buffer[84]) );
  DFFRX1 out_buffer_reg_10__5_ ( .D(N632), .CK(GCK), .RN(n408), .Q(
        out_buffer[85]) );
  DFFRX1 out_buffer_reg_10__7_ ( .D(N634), .CK(GCK), .RN(n408), .Q(
        out_buffer[87]) );
  DFFRX1 out_buffer_reg_9__4_ ( .D(N581), .CK(GCK), .RN(n4100), .Q(
        out_buffer[100]) );
  DFFRX1 out_buffer_reg_8__4_ ( .D(N531), .CK(GCK), .RN(n4110), .Q(
        out_buffer[116]) );
  DFFRX1 out_buffer_reg_8__5_ ( .D(N532), .CK(GCK), .RN(n4110), .Q(
        out_buffer[117]) );
  DFFRX1 out_buffer_reg_8__7_ ( .D(N534), .CK(GCK), .RN(n4110), .Q(
        out_buffer[119]) );
  DFFRX1 out_buffer_reg_8__9_ ( .D(N536), .CK(GCK), .RN(n4110), .Q(
        out_buffer[121]) );
  DFFRX1 out_buffer_reg_7__4_ ( .D(N481), .CK(GCK), .RN(n4120), .Q(
        out_buffer[132]) );
  DFFRX1 out_buffer_reg_7__5_ ( .D(N482), .CK(GCK), .RN(n4130), .Q(
        out_buffer[133]) );
  DFFRX1 out_buffer_reg_7__7_ ( .D(N484), .CK(GCK), .RN(n4130), .Q(
        out_buffer[135]) );
  DFFRX1 out_buffer_reg_7__9_ ( .D(N486), .CK(GCK), .RN(n4130), .Q(
        out_buffer[137]) );
  DFFRX1 out_buffer_reg_6__4_ ( .D(N431), .CK(GCK), .RN(n4140), .Q(
        out_buffer[148]) );
  DFFRX1 out_buffer_reg_6__5_ ( .D(N432), .CK(GCK), .RN(n4140), .Q(
        out_buffer[149]) );
  DFFRX1 out_buffer_reg_6__6_ ( .D(N433), .CK(GCK), .RN(n4140), .Q(
        out_buffer[150]) );
  DFFRX1 out_buffer_reg_5__4_ ( .D(N381), .CK(GCK), .RN(n4150), .Q(
        out_buffer[164]) );
  DFFRX1 out_buffer_reg_5__6_ ( .D(N383), .CK(GCK), .RN(n4150), .Q(
        out_buffer[166]) );
  DFFRX1 out_buffer_reg_4__7_ ( .D(N334), .CK(GCK), .RN(n4170), .Q(
        out_buffer[183]) );
  DFFRX1 out_buffer_reg_3__4_ ( .D(N281), .CK(GCK), .RN(n4180), .Q(
        out_buffer[196]) );
  DFFRX1 out_buffer_reg_3__5_ ( .D(N282), .CK(GCK), .RN(n4180), .Q(
        out_buffer[197]) );
  DFFRX1 out_buffer_reg_3__7_ ( .D(N284), .CK(GCK), .RN(n4180), .Q(
        out_buffer[199]) );
  DFFRX1 out_buffer_reg_3__9_ ( .D(N286), .CK(GCK), .RN(n4190), .Q(
        out_buffer[201]) );
  DFFRX1 out_buffer_reg_2__4_ ( .D(N231), .CK(GCK), .RN(n4200), .Q(
        out_buffer[212]) );
  DFFRX1 out_buffer_reg_2__5_ ( .D(N232), .CK(GCK), .RN(n4200), .Q(
        out_buffer[213]) );
  DFFRX1 out_buffer_reg_2__7_ ( .D(N234), .CK(GCK), .RN(n4200), .Q(
        out_buffer[215]) );
  DFFRX1 out_buffer_reg_2__9_ ( .D(N236), .CK(GCK), .RN(n4200), .Q(
        out_buffer[217]) );
  DFFRX1 out_buffer_reg_1__5_ ( .D(N182), .CK(GCK), .RN(n4210), .Q(
        out_buffer[229]) );
  DFFRX1 out_buffer_reg_1__7_ ( .D(N184), .CK(GCK), .RN(n4210), .Q(
        out_buffer[231]) );
  DFFRX1 out_buffer_reg_1__9_ ( .D(N186), .CK(GCK), .RN(n4210), .Q(
        out_buffer[233]) );
  DFFRX1 out_buffer_reg_0__4_ ( .D(N131), .CK(GCK), .RN(n4220), .Q(
        out_buffer[244]) );
  DFFRX1 out_buffer_reg_0__5_ ( .D(N132), .CK(GCK), .RN(n4220), .Q(
        out_buffer[245]) );
  DFFRX1 out_buffer_reg_0__7_ ( .D(N134), .CK(GCK), .RN(n4230), .Q(
        out_buffer[247]) );
  DFFRX1 out_buffer_reg_0__9_ ( .D(N136), .CK(GCK), .RN(n4230), .Q(
        out_buffer[249]) );
  DFFRX1 rd_addr_reg_2_ ( .D(n1089), .CK(GCK), .RN(n400), .Q(addr[2]), .QN(n6)
         );
  DFFRX1 rd_addr_reg_3_ ( .D(n1088), .CK(GCK), .RN(n400), .Q(addr[3]), .QN(n7)
         );
  DFFRX1 out_buffer_reg_13__3_ ( .D(N780), .CK(GCK), .RN(n404), .Q(
        out_buffer[35]) );
  DFFRX1 out_buffer_reg_11__3_ ( .D(N680), .CK(GCK), .RN(n407), .Q(
        out_buffer[67]) );
  DFFRX1 out_buffer_reg_10__2_ ( .D(N629), .CK(GCK), .RN(n408), .Q(
        out_buffer[82]) );
  DFFRX1 out_buffer_reg_9__3_ ( .D(N580), .CK(GCK), .RN(n4100), .Q(
        out_buffer[99]) );
  DFFRX1 out_buffer_reg_8__3_ ( .D(N530), .CK(GCK), .RN(n4110), .Q(
        out_buffer[115]) );
  DFFRX1 out_buffer_reg_7__1_ ( .D(N478), .CK(GCK), .RN(n4120), .Q(
        out_buffer[129]) );
  DFFRX1 out_buffer_reg_7__3_ ( .D(N480), .CK(GCK), .RN(n4120), .Q(
        out_buffer[131]) );
  DFFRX1 out_buffer_reg_6__3_ ( .D(N430), .CK(GCK), .RN(n4140), .Q(
        out_buffer[147]) );
  DFFRX1 out_buffer_reg_4__3_ ( .D(N330), .CK(GCK), .RN(n4170), .Q(
        out_buffer[179]) );
  DFFRX1 out_buffer_reg_3__3_ ( .D(N280), .CK(GCK), .RN(n4180), .Q(
        out_buffer[195]) );
  DFFRX1 out_buffer_reg_2__1_ ( .D(N228), .CK(GCK), .RN(n4190), .Q(
        out_buffer[209]) );
  DFFRX1 out_buffer_reg_2__3_ ( .D(N230), .CK(GCK), .RN(n4190), .Q(
        out_buffer[211]) );
  DFFRX1 out_buffer_reg_1__3_ ( .D(N180), .CK(GCK), .RN(n4210), .Q(
        out_buffer[227]) );
  DFFRX1 out_buffer_reg_0__3_ ( .D(N130), .CK(GCK), .RN(n4220), .Q(
        out_buffer[243]) );
  DFFRX1 out_buffer_reg_15__0_ ( .D(N877), .CK(GCK), .RN(n401), .Q(
        out_buffer[0]) );
  DFFRX1 out_buffer_reg_13__0_ ( .D(N777), .CK(GCK), .RN(n404), .Q(
        out_buffer[32]) );
  DFFRX1 out_buffer_reg_11__0_ ( .D(N677), .CK(GCK), .RN(n406), .Q(
        out_buffer[64]) );
  DFFRX1 out_buffer_reg_8__0_ ( .D(N527), .CK(GCK), .RN(n4110), .Q(
        out_buffer[112]) );
  DFFRX1 out_buffer_reg_7__0_ ( .D(N477), .CK(GCK), .RN(n4120), .Q(
        out_buffer[128]) );
  DFFRX1 out_buffer_reg_3__0_ ( .D(N277), .CK(GCK), .RN(n4180), .Q(
        out_buffer[192]) );
  DFFRX1 out_buffer_reg_2__0_ ( .D(N227), .CK(GCK), .RN(n4190), .Q(
        out_buffer[208]) );
  DFFRX1 out_buffer_reg_1__0_ ( .D(N177), .CK(GCK), .RN(n4210), .Q(
        out_buffer[224]) );
  DFFRX1 out_cs_reg_2_ ( .D(n1093), .CK(GCK), .RN(n399), .Q(out_cs[2]), .QN(
        n96) );
  DFFRX1 out_cs_reg_1_ ( .D(n1092), .CK(GCK), .RN(n399), .Q(out_cs[1]), .QN(
        n88) );
  DFFRX1 out_buffer_reg_10__13_ ( .D(N640), .CK(GCK), .RN(n409), .Q(
        out_buffer[93]) );
  DFFRX1 out_buffer_reg_9__13_ ( .D(N590), .CK(GCK), .RN(n4100), .Q(
        out_buffer[109]) );
  DFFRX1 out_buffer_reg_6__13_ ( .D(N440), .CK(GCK), .RN(n4150), .Q(
        out_buffer[157]) );
  DFFRX1 out_buffer_reg_5__13_ ( .D(N390), .CK(GCK), .RN(n4160), .Q(
        out_buffer[173]) );
  DFFRX1 out_buffer_reg_14__13_ ( .D(N840), .CK(GCK), .RN(n403), .Q(
        out_buffer[29]) );
  DFFRX1 out_buffer_reg_12__3_ ( .D(N730), .CK(GCK), .RN(n405), .Q(
        out_buffer[51]) );
  DFFRX1 out_buffer_reg_10__3_ ( .D(N630), .CK(GCK), .RN(n408), .Q(
        out_buffer[83]) );
  DFFRX1 out_buffer_reg_6__2_ ( .D(N429), .CK(GCK), .RN(n4140), .Q(
        out_buffer[146]) );
  DFFRX1 out_buffer_reg_5__2_ ( .D(N379), .CK(GCK), .RN(n4150), .Q(
        out_buffer[162]) );
  DFFRX1 out_buffer_reg_14__2_ ( .D(N829), .CK(GCK), .RN(n402), .Q(
        out_buffer[18]) );
  DFFRX1 out_buffer_reg_6__8_ ( .D(N435), .CK(GCK), .RN(n4140), .Q(
        out_buffer[152]) );
  DFFRX1 out_buffer_reg_5__8_ ( .D(N385), .CK(GCK), .RN(n4160), .Q(
        out_buffer[168]) );
  DFFRX1 out_buffer_reg_6__11_ ( .D(N438), .CK(GCK), .RN(n4140), .Q(
        out_buffer[155]) );
  DFFRX1 out_buffer_reg_5__11_ ( .D(N388), .CK(GCK), .RN(n4160), .Q(
        out_buffer[171]) );
  DFFRX1 out_buffer_reg_14__4_ ( .D(N831), .CK(GCK), .RN(n403), .Q(
        out_buffer[20]) );
  DFFRX1 out_buffer_reg_14__8_ ( .D(N835), .CK(GCK), .RN(n403), .Q(
        out_buffer[24]) );
  DFFRX1 out_buffer_reg_14__15_ ( .D(N842), .CK(GCK), .RN(n403), .Q(
        out_buffer[31]) );
  DFFRX1 out_buffer_reg_12__12_ ( .D(N739), .CK(GCK), .RN(n406), .Q(
        out_buffer[60]) );
  DFFRX1 out_buffer_reg_10__12_ ( .D(N639), .CK(GCK), .RN(n409), .Q(
        out_buffer[92]) );
  DFFRX1 out_buffer_reg_14__9_ ( .D(N836), .CK(GCK), .RN(n403), .Q(
        out_buffer[25]) );
  DFFRX1 out_buffer_reg_5__15_ ( .D(N392), .CK(GCK), .RN(n4160), .Q(
        out_buffer[175]) );
  DFFRX1 out_buffer_reg_5__9_ ( .D(N386), .CK(GCK), .RN(n4160), .Q(
        out_buffer[169]) );
  DFFRX1 out_buffer_reg_14__3_ ( .D(N830), .CK(GCK), .RN(n402), .Q(
        out_buffer[19]) );
  DFFRX1 out_buffer_reg_6__7_ ( .D(N434), .CK(GCK), .RN(n4140), .Q(
        out_buffer[151]) );
  DFFRX1 out_buffer_reg_5__7_ ( .D(N384), .CK(GCK), .RN(n4160), .Q(
        out_buffer[167]) );
  DFFRX1 out_buffer_reg_6__9_ ( .D(N436), .CK(GCK), .RN(n4140), .Q(
        out_buffer[153]) );
  DFFRX1 out_buffer_reg_6__10_ ( .D(N437), .CK(GCK), .RN(n4140), .Q(
        out_buffer[154]) );
  DFFRX1 out_buffer_reg_14__11_ ( .D(N838), .CK(GCK), .RN(n403), .Q(
        out_buffer[27]) );
  DFFRX1 out_buffer_reg_5__3_ ( .D(N380), .CK(GCK), .RN(n4150), .Q(
        out_buffer[163]) );
  DFFRX1 out_buffer_reg_14__6_ ( .D(N833), .CK(GCK), .RN(n403), .Q(
        out_buffer[22]) );
  DFFRX1 out_buffer_reg_12__8_ ( .D(N735), .CK(GCK), .RN(n406), .Q(
        out_buffer[56]) );
  DFFRX1 out_buffer_reg_14__10_ ( .D(N837), .CK(GCK), .RN(n403), .Q(
        out_buffer[26]) );
  DFFRX1 out_buffer_reg_9__7_ ( .D(N584), .CK(GCK), .RN(n4100), .Q(
        out_buffer[103]) );
  DFFRX1 out_buffer_reg_5__5_ ( .D(N382), .CK(GCK), .RN(n4150), .Q(
        out_buffer[165]) );
  DFFRX1 out_buffer_reg_10__8_ ( .D(N635), .CK(GCK), .RN(n409), .Q(
        out_buffer[88]) );
  DFFRX1 out_buffer_reg_9__11_ ( .D(N588), .CK(GCK), .RN(n4100), .Q(
        out_buffer[107]) );
  DFFRX1 out_buffer_reg_9__6_ ( .D(N583), .CK(GCK), .RN(n4100), .Q(
        out_buffer[102]) );
  DFFRX1 out_buffer_reg_9__9_ ( .D(N586), .CK(GCK), .RN(n4100), .Q(
        out_buffer[105]) );
  DFFRX1 out_buffer_reg_10__9_ ( .D(N636), .CK(GCK), .RN(n409), .Q(
        out_buffer[89]) );
  DFFRX1 out_buffer_reg_10__15_ ( .D(N642), .CK(GCK), .RN(n409), .Q(
        out_buffer[95]) );
  DFFRX1 out_buffer_reg_6__15_ ( .D(N442), .CK(GCK), .RN(n4150), .Q(
        out_buffer[159]) );
  DFFRX1 out_buffer_reg_14__12_ ( .D(N839), .CK(GCK), .RN(n403), .Q(
        out_buffer[28]) );
  DFFRX1 out_buffer_reg_9__10_ ( .D(N587), .CK(GCK), .RN(n4100), .Q(
        out_buffer[106]) );
  DFFRX1 out_buffer_reg_5__10_ ( .D(N387), .CK(GCK), .RN(n4160), .Q(
        out_buffer[170]) );
  DFFRX2 rd_addr_reg_0_ ( .D(n1091), .CK(GCK), .RN(n399), .Q(addr[0]), .QN(n4)
         );
  DFFRX2 rd_addr_reg_10_ ( .D(n1081), .CK(GCK), .RN(n400), .Q(rd_addr[10]) );
  DFFRX2 rd_reg_reg_15__15_ ( .D(n1067), .CK(GCK), .RN(n400), .QN(n5890) );
  DFFRX2 rd_addr_reg_1_ ( .D(n1090), .CK(GCK), .RN(n399), .Q(addr[1]), .QN(n5)
         );
  DFFRX1 en_reg ( .D(N45), .CK(GCK), .RN(n109), .Q(en) );
  DFFRX1 cnt_reg_0_ ( .D(N39), .CK(GCK), .RN(n108), .Q(cnt[0]) );
  DFFRX1 r_push_buffer_reg ( .D(n1075), .CK(GCK), .RN(n107), .Q(n90), .QN(
        n5880) );
  DFFRX1 cnt_reg_1_ ( .D(N40), .CK(GCK), .RN(n109), .Q(cnt[1]) );
  DFFRX1 cnt_reg_2_ ( .D(N41), .CK(GCK), .RN(n108), .Q(cnt[2]) );
  DFFRX1 rd_reg_reg_14__6_ ( .D(n922), .CK(GCK), .RN(n107), .Q(rd_reg[21]), 
        .QN(n7160) );
  DFFRX1 rd_reg_reg_14__5_ ( .D(n906), .CK(GCK), .RN(n109), .Q(rd_reg[20]), 
        .QN(n7300) );
  DFFRX1 rd_reg_reg_13__5_ ( .D(n905), .CK(GCK), .RN(n108), .Q(rd_reg[36]), 
        .QN(n7310) );
  DFFRX1 rd_reg_reg_12__6_ ( .D(n920), .CK(GCK), .RN(n107), .Q(rd_reg[53]), 
        .QN(n7180) );
  DFFRX1 rd_reg_reg_12__5_ ( .D(n904), .CK(GCK), .RN(n109), .Q(rd_reg[52]), 
        .QN(n7320) );
  DFFRX1 rd_reg_reg_11__5_ ( .D(n903), .CK(GCK), .RN(n108), .Q(rd_reg[68]), 
        .QN(n7330) );
  DFFRX1 rd_reg_reg_9__6_ ( .D(n917), .CK(GCK), .RN(n107), .Q(rd_reg[101]), 
        .QN(n7210) );
  DFFRX1 rd_reg_reg_6__6_ ( .D(n914), .CK(GCK), .RN(n109), .Q(rd_reg[149]), 
        .QN(n7240) );
  DFFRX1 rd_reg_reg_5__6_ ( .D(n913), .CK(GCK), .RN(n108), .Q(rd_reg[165]), 
        .QN(n7250) );
  DFFRX1 rd_reg_reg_3__6_ ( .D(n911), .CK(GCK), .RN(n107), .Q(rd_reg[197]), 
        .QN(n7270) );
  DFFRX1 rd_reg_reg_2__7_ ( .D(n926), .CK(GCK), .RN(n109), .Q(rd_reg[214]), 
        .QN(n7140) );
  DFFRX1 rd_reg_reg_2__6_ ( .D(n910), .CK(GCK), .RN(n108), .Q(rd_reg[213]), 
        .QN(n7280) );
  DFFRX1 rd_reg_reg_1__6_ ( .D(n909), .CK(GCK), .RN(n107), .Q(rd_reg[229]), 
        .QN(n7290) );
  DFFRX1 rd_reg_reg_0__12_ ( .D(n1004), .CK(GCK), .RN(n109), .Q(rd_reg[251])
         );
  DFFRX1 rd_reg_reg_0__11_ ( .D(n988), .CK(GCK), .RN(n108), .Q(rd_reg[250]) );
  DFFRX1 rd_reg_reg_0__10_ ( .D(n972), .CK(GCK), .RN(n107), .Q(rd_reg[249]) );
  DFFRX1 rd_reg_reg_0__14_ ( .D(n1036), .CK(GCK), .RN(n109), .Q(rd_reg[253])
         );
  DFFRX1 rd_reg_reg_0__2_ ( .D(n844), .CK(GCK), .RN(n108), .Q(rd_reg[241]) );
  DFFRX1 rd_reg_reg_0__1_ ( .D(n8280), .CK(GCK), .RN(n107), .Q(rd_reg[240]) );
  DFFRX1 rd_reg_reg_0__15_ ( .D(n1052), .CK(GCK), .RN(n109), .Q(rd_reg[254])
         );
  DFFRX1 rd_reg_reg_0__13_ ( .D(n1020), .CK(GCK), .RN(n108), .Q(rd_reg[252])
         );
  DFFRX1 rd_reg_reg_0__9_ ( .D(n956), .CK(GCK), .RN(n107), .Q(rd_reg[248]) );
  DFFRX1 rd_reg_reg_0__8_ ( .D(n940), .CK(GCK), .RN(n109), .Q(rd_reg[247]) );
  DFFRX1 rd_reg_reg_0__7_ ( .D(n924), .CK(GCK), .RN(n108), .Q(rd_reg[246]) );
  DFFRX1 rd_reg_reg_0__6_ ( .D(n908), .CK(GCK), .RN(n107), .Q(rd_reg[245]) );
  DFFRX1 rd_reg_reg_0__5_ ( .D(n8920), .CK(GCK), .RN(n109), .Q(rd_reg[244]) );
  DFFRX1 rd_reg_reg_0__4_ ( .D(n8760), .CK(GCK), .RN(n108), .Q(rd_reg[243]) );
  DFFRX1 rd_reg_reg_0__3_ ( .D(n8600), .CK(GCK), .RN(n107), .Q(rd_reg[242]) );
  DFFRX1 rd_reg_reg_0__0_ ( .D(n8120), .CK(GCK), .RN(n109), .Q(rd_reg[239]) );
  DFFRX1 rd_reg_reg_13__6_ ( .D(n921), .CK(GCK), .RN(n108), .Q(rd_reg[37]), 
        .QN(n7170) );
  DFFRX1 rd_reg_reg_11__6_ ( .D(n919), .CK(GCK), .RN(n107), .Q(rd_reg[69]), 
        .QN(n7190) );
  DFFRX1 rd_reg_reg_10__6_ ( .D(n918), .CK(GCK), .RN(n109), .Q(rd_reg[85]), 
        .QN(n7200) );
  DFFRX1 rd_reg_reg_8__6_ ( .D(n916), .CK(GCK), .RN(n108), .Q(rd_reg[117]), 
        .QN(n7220) );
  DFFRX1 rd_reg_reg_4__6_ ( .D(n912), .CK(GCK), .RN(n107), .Q(rd_reg[181]), 
        .QN(n7260) );
  DFFRX1 rd_reg_reg_3__7_ ( .D(n927), .CK(GCK), .RN(n109), .Q(rd_reg[198]), 
        .QN(n7130) );
  DFFRX1 rd_reg_reg_1__7_ ( .D(n925), .CK(GCK), .RN(n108), .Q(rd_reg[230]), 
        .QN(n7150) );
  DFFRX1 rd_reg_reg_14__14_ ( .D(n1050), .CK(GCK), .RN(n107), .Q(rd_reg[29]), 
        .QN(n604) );
  DFFRX1 rd_reg_reg_14__13_ ( .D(n1034), .CK(GCK), .RN(n109), .Q(rd_reg[28]), 
        .QN(n6180) );
  DFFRX1 rd_reg_reg_14__12_ ( .D(n1018), .CK(GCK), .RN(n108), .Q(rd_reg[27]), 
        .QN(n6320) );
  DFFRX1 rd_reg_reg_14__11_ ( .D(n1002), .CK(GCK), .RN(n107), .Q(rd_reg[26]), 
        .QN(n646) );
  DFFRX1 rd_reg_reg_14__10_ ( .D(n986), .CK(GCK), .RN(n109), .Q(rd_reg[25]), 
        .QN(n6600) );
  DFFRX1 rd_reg_reg_14__9_ ( .D(n970), .CK(GCK), .RN(n108), .Q(rd_reg[24]), 
        .QN(n6740) );
  DFFRX1 rd_reg_reg_14__8_ ( .D(n954), .CK(GCK), .RN(n107), .Q(rd_reg[23]), 
        .QN(n6880) );
  DFFRX1 rd_reg_reg_14__7_ ( .D(n938), .CK(GCK), .RN(n109), .Q(rd_reg[22]), 
        .QN(n702) );
  DFFRX1 rd_reg_reg_14__1_ ( .D(n8420), .CK(GCK), .RN(n108), .Q(rd_reg[16]), 
        .QN(n7860) );
  DFFRX1 rd_reg_reg_13__14_ ( .D(n1049), .CK(GCK), .RN(n107), .Q(rd_reg[45]), 
        .QN(n605) );
  DFFRX1 rd_reg_reg_13__13_ ( .D(n1033), .CK(GCK), .RN(n109), .Q(rd_reg[44]), 
        .QN(n6190) );
  DFFRX1 rd_reg_reg_13__12_ ( .D(n1017), .CK(GCK), .RN(n108), .Q(rd_reg[43]), 
        .QN(n6330) );
  DFFRX1 rd_reg_reg_13__11_ ( .D(n1001), .CK(GCK), .RN(n107), .Q(rd_reg[42]), 
        .QN(n647) );
  DFFRX1 rd_reg_reg_13__10_ ( .D(n985), .CK(GCK), .RN(n109), .Q(rd_reg[41]), 
        .QN(n6610) );
  DFFRX1 rd_reg_reg_13__9_ ( .D(n969), .CK(GCK), .RN(n108), .Q(rd_reg[40]), 
        .QN(n6750) );
  DFFRX1 rd_reg_reg_13__8_ ( .D(n953), .CK(GCK), .RN(n107), .Q(rd_reg[39]), 
        .QN(n6890) );
  DFFRX1 rd_reg_reg_13__7_ ( .D(n937), .CK(GCK), .RN(n109), .Q(rd_reg[38]), 
        .QN(n703) );
  DFFRX1 rd_reg_reg_13__1_ ( .D(n8410), .CK(GCK), .RN(n108), .Q(rd_reg[32]), 
        .QN(n7870) );
  DFFRX1 rd_reg_reg_12__14_ ( .D(n1048), .CK(GCK), .RN(n107), .Q(rd_reg[61]), 
        .QN(n606) );
  DFFRX1 rd_reg_reg_12__13_ ( .D(n1032), .CK(GCK), .RN(n109), .Q(rd_reg[60]), 
        .QN(n6200) );
  DFFRX1 rd_reg_reg_12__12_ ( .D(n1016), .CK(GCK), .RN(n108), .Q(rd_reg[59]), 
        .QN(n6340) );
  DFFRX1 rd_reg_reg_12__11_ ( .D(n1000), .CK(GCK), .RN(n107), .Q(rd_reg[58]), 
        .QN(n648) );
  DFFRX1 rd_reg_reg_12__10_ ( .D(n984), .CK(GCK), .RN(n109), .Q(rd_reg[57]), 
        .QN(n6620) );
  DFFRX1 rd_reg_reg_12__9_ ( .D(n968), .CK(GCK), .RN(n108), .Q(rd_reg[56]), 
        .QN(n6760) );
  DFFRX1 rd_reg_reg_12__8_ ( .D(n952), .CK(GCK), .RN(n107), .Q(rd_reg[55]), 
        .QN(n6900) );
  DFFRX1 rd_reg_reg_12__7_ ( .D(n936), .CK(GCK), .RN(n109), .Q(rd_reg[54]), 
        .QN(n704) );
  DFFRX1 rd_reg_reg_12__1_ ( .D(n8400), .CK(GCK), .RN(n108), .Q(rd_reg[48]), 
        .QN(n7880) );
  DFFRX1 rd_reg_reg_12__0_ ( .D(n8240), .CK(GCK), .RN(n107), .Q(rd_reg[47]), 
        .QN(n801) );
  DFFRX1 rd_reg_reg_11__14_ ( .D(n1047), .CK(GCK), .RN(n109), .Q(rd_reg[77]), 
        .QN(n607) );
  DFFRX1 rd_reg_reg_11__13_ ( .D(n1031), .CK(GCK), .RN(n108), .Q(rd_reg[76]), 
        .QN(n6210) );
  DFFRX1 rd_reg_reg_11__12_ ( .D(n1015), .CK(GCK), .RN(n107), .Q(rd_reg[75]), 
        .QN(n6350) );
  DFFRX1 rd_reg_reg_11__11_ ( .D(n999), .CK(GCK), .RN(n109), .Q(rd_reg[74]), 
        .QN(n649) );
  DFFRX1 rd_reg_reg_11__10_ ( .D(n983), .CK(GCK), .RN(n108), .Q(rd_reg[73]), 
        .QN(n6630) );
  DFFRX1 rd_reg_reg_11__9_ ( .D(n967), .CK(GCK), .RN(n107), .Q(rd_reg[72]), 
        .QN(n6770) );
  DFFRX1 rd_reg_reg_11__8_ ( .D(n951), .CK(GCK), .RN(n109), .Q(rd_reg[71]), 
        .QN(n6910) );
  DFFRX1 rd_reg_reg_11__1_ ( .D(n8390), .CK(GCK), .RN(n108), .Q(rd_reg[64]), 
        .QN(n7890) );
  DFFRX1 rd_reg_reg_11__0_ ( .D(n8230), .CK(GCK), .RN(n107), .Q(rd_reg[63]), 
        .QN(n802) );
  DFFRX1 rd_reg_reg_10__14_ ( .D(n1046), .CK(GCK), .RN(n109), .Q(rd_reg[93]), 
        .QN(n608) );
  DFFRX1 rd_reg_reg_10__13_ ( .D(n1030), .CK(GCK), .RN(n108), .Q(rd_reg[92]), 
        .QN(n6220) );
  DFFRX1 rd_reg_reg_10__12_ ( .D(n1014), .CK(GCK), .RN(n107), .Q(rd_reg[91]), 
        .QN(n6360) );
  DFFRX1 rd_reg_reg_10__11_ ( .D(n998), .CK(GCK), .RN(n109), .Q(rd_reg[90]), 
        .QN(n650) );
  DFFRX1 rd_reg_reg_10__10_ ( .D(n982), .CK(GCK), .RN(n108), .Q(rd_reg[89]), 
        .QN(n6640) );
  DFFRX1 rd_reg_reg_10__9_ ( .D(n966), .CK(GCK), .RN(n107), .Q(rd_reg[88]), 
        .QN(n6780) );
  DFFRX1 rd_reg_reg_10__8_ ( .D(n950), .CK(GCK), .RN(n109), .Q(rd_reg[87]), 
        .QN(n6920) );
  DFFRX1 rd_reg_reg_10__1_ ( .D(n8380), .CK(GCK), .RN(n108), .Q(rd_reg[80]), 
        .QN(n7900) );
  DFFRX1 rd_reg_reg_10__0_ ( .D(n8220), .CK(GCK), .RN(n107), .Q(rd_reg[79]), 
        .QN(n803) );
  DFFRX1 rd_reg_reg_9__14_ ( .D(n1045), .CK(GCK), .RN(n109), .Q(rd_reg[109]), 
        .QN(n609) );
  DFFRX1 rd_reg_reg_9__13_ ( .D(n1029), .CK(GCK), .RN(n108), .Q(rd_reg[108]), 
        .QN(n6230) );
  DFFRX1 rd_reg_reg_9__12_ ( .D(n1013), .CK(GCK), .RN(n107), .Q(rd_reg[107]), 
        .QN(n6370) );
  DFFRX1 rd_reg_reg_9__11_ ( .D(n997), .CK(GCK), .RN(n109), .Q(rd_reg[106]), 
        .QN(n651) );
  DFFRX1 rd_reg_reg_9__10_ ( .D(n981), .CK(GCK), .RN(n108), .Q(rd_reg[105]), 
        .QN(n6650) );
  DFFRX1 rd_reg_reg_9__9_ ( .D(n965), .CK(GCK), .RN(n107), .Q(rd_reg[104]), 
        .QN(n6790) );
  DFFRX1 rd_reg_reg_9__8_ ( .D(n949), .CK(GCK), .RN(n109), .Q(rd_reg[103]), 
        .QN(n6930) );
  DFFRX1 rd_reg_reg_9__1_ ( .D(n8370), .CK(GCK), .RN(n108), .Q(rd_reg[96]), 
        .QN(n7910) );
  DFFRX1 rd_reg_reg_9__0_ ( .D(n8210), .CK(GCK), .RN(n107), .Q(rd_reg[95]), 
        .QN(n804) );
  DFFRX1 rd_reg_reg_8__14_ ( .D(n1044), .CK(GCK), .RN(n109), .Q(rd_reg[125]), 
        .QN(n6100) );
  DFFRX1 rd_reg_reg_8__13_ ( .D(n1028), .CK(GCK), .RN(n108), .Q(rd_reg[124]), 
        .QN(n6240) );
  DFFRX1 rd_reg_reg_8__12_ ( .D(n1012), .CK(GCK), .RN(n107), .Q(rd_reg[123]), 
        .QN(n6380) );
  DFFRX1 rd_reg_reg_8__11_ ( .D(n996), .CK(GCK), .RN(n109), .Q(rd_reg[122]), 
        .QN(n652) );
  DFFRX1 rd_reg_reg_8__10_ ( .D(n980), .CK(GCK), .RN(n108), .Q(rd_reg[121]), 
        .QN(n6660) );
  DFFRX1 rd_reg_reg_8__9_ ( .D(n964), .CK(GCK), .RN(n107), .Q(rd_reg[120]), 
        .QN(n6800) );
  DFFRX1 rd_reg_reg_8__8_ ( .D(n948), .CK(GCK), .RN(n109), .Q(rd_reg[119]), 
        .QN(n694) );
  DFFRX1 rd_reg_reg_8__1_ ( .D(n8360), .CK(GCK), .RN(n108), .Q(rd_reg[112]), 
        .QN(n7920) );
  DFFRX1 rd_reg_reg_8__0_ ( .D(n8200), .CK(GCK), .RN(n107), .Q(rd_reg[111]), 
        .QN(n805) );
  DFFRX1 rd_reg_reg_7__14_ ( .D(n1043), .CK(GCK), .RN(n109), .Q(rd_reg[141]), 
        .QN(n6110) );
  DFFRX1 rd_reg_reg_7__13_ ( .D(n1027), .CK(GCK), .RN(n108), .Q(rd_reg[140]), 
        .QN(n6250) );
  DFFRX1 rd_reg_reg_7__12_ ( .D(n1011), .CK(GCK), .RN(n107), .Q(rd_reg[139]), 
        .QN(n6390) );
  DFFRX1 rd_reg_reg_7__11_ ( .D(n995), .CK(GCK), .RN(n109), .Q(rd_reg[138]), 
        .QN(n653) );
  DFFRX1 rd_reg_reg_7__10_ ( .D(n979), .CK(GCK), .RN(n108), .Q(rd_reg[137]), 
        .QN(n6670) );
  DFFRX1 rd_reg_reg_7__9_ ( .D(n963), .CK(GCK), .RN(n107), .Q(rd_reg[136]), 
        .QN(n6810) );
  DFFRX1 rd_reg_reg_7__8_ ( .D(n947), .CK(GCK), .RN(n109), .Q(rd_reg[135]), 
        .QN(n695) );
  DFFRX1 rd_reg_reg_7__1_ ( .D(n8350), .CK(GCK), .RN(n108), .Q(rd_reg[128]), 
        .QN(n7930) );
  DFFRX1 rd_reg_reg_7__0_ ( .D(n8190), .CK(GCK), .RN(n107), .Q(rd_reg[127]), 
        .QN(n806) );
  DFFRX1 rd_reg_reg_6__14_ ( .D(n1042), .CK(GCK), .RN(n109), .Q(rd_reg[157]), 
        .QN(n6120) );
  DFFRX1 rd_reg_reg_6__13_ ( .D(n1026), .CK(GCK), .RN(n108), .Q(rd_reg[156]), 
        .QN(n6260) );
  DFFRX1 rd_reg_reg_6__12_ ( .D(n1010), .CK(GCK), .RN(n107), .Q(rd_reg[155]), 
        .QN(n6400) );
  DFFRX1 rd_reg_reg_6__11_ ( .D(n994), .CK(GCK), .RN(n109), .Q(rd_reg[154]), 
        .QN(n654) );
  DFFRX1 rd_reg_reg_6__10_ ( .D(n978), .CK(GCK), .RN(n108), .Q(rd_reg[153]), 
        .QN(n6680) );
  DFFRX1 rd_reg_reg_6__9_ ( .D(n962), .CK(GCK), .RN(n107), .Q(rd_reg[152]), 
        .QN(n6820) );
  DFFRX1 rd_reg_reg_6__8_ ( .D(n946), .CK(GCK), .RN(n109), .Q(rd_reg[151]), 
        .QN(n696) );
  DFFRX1 rd_reg_reg_6__1_ ( .D(n8340), .CK(GCK), .RN(n108), .Q(rd_reg[144]), 
        .QN(n794) );
  DFFRX1 rd_reg_reg_6__0_ ( .D(n8180), .CK(GCK), .RN(n107), .Q(rd_reg[143]), 
        .QN(n807) );
  DFFRX1 rd_reg_reg_5__14_ ( .D(n1041), .CK(GCK), .RN(n109), .Q(rd_reg[173]), 
        .QN(n6130) );
  DFFRX1 rd_reg_reg_5__13_ ( .D(n1025), .CK(GCK), .RN(n108), .Q(rd_reg[172]), 
        .QN(n6270) );
  DFFRX1 rd_reg_reg_5__12_ ( .D(n1009), .CK(GCK), .RN(n107), .Q(rd_reg[171]), 
        .QN(n6410) );
  DFFRX1 rd_reg_reg_5__11_ ( .D(n993), .CK(GCK), .RN(n109), .Q(rd_reg[170]), 
        .QN(n655) );
  DFFRX1 rd_reg_reg_5__10_ ( .D(n977), .CK(GCK), .RN(n108), .Q(rd_reg[169]), 
        .QN(n6690) );
  DFFRX1 rd_reg_reg_5__9_ ( .D(n961), .CK(GCK), .RN(n107), .Q(rd_reg[168]), 
        .QN(n6830) );
  DFFRX1 rd_reg_reg_5__8_ ( .D(n945), .CK(GCK), .RN(n109), .Q(rd_reg[167]), 
        .QN(n697) );
  DFFRX1 rd_reg_reg_5__7_ ( .D(n929), .CK(GCK), .RN(n108), .Q(rd_reg[166]), 
        .QN(n7110) );
  DFFRX1 rd_reg_reg_5__1_ ( .D(n8330), .CK(GCK), .RN(n107), .Q(rd_reg[160]), 
        .QN(n795) );
  DFFRX1 rd_reg_reg_5__0_ ( .D(n8170), .CK(GCK), .RN(n109), .Q(rd_reg[159]), 
        .QN(n808) );
  DFFRX1 rd_reg_reg_4__14_ ( .D(n1040), .CK(GCK), .RN(n108), .Q(rd_reg[189]), 
        .QN(n6140) );
  DFFRX1 rd_reg_reg_4__13_ ( .D(n1024), .CK(GCK), .RN(n107), .Q(rd_reg[188]), 
        .QN(n6280) );
  DFFRX1 rd_reg_reg_4__12_ ( .D(n1008), .CK(GCK), .RN(n109), .Q(rd_reg[187]), 
        .QN(n6420) );
  DFFRX1 rd_reg_reg_4__11_ ( .D(n992), .CK(GCK), .RN(n108), .Q(rd_reg[186]), 
        .QN(n656) );
  DFFRX1 rd_reg_reg_4__10_ ( .D(n976), .CK(GCK), .RN(n107), .Q(rd_reg[185]), 
        .QN(n6700) );
  DFFRX1 rd_reg_reg_4__9_ ( .D(n960), .CK(GCK), .RN(n109), .Q(rd_reg[184]), 
        .QN(n6840) );
  DFFRX1 rd_reg_reg_4__8_ ( .D(n944), .CK(GCK), .RN(n108), .Q(rd_reg[183]), 
        .QN(n698) );
  DFFRX1 rd_reg_reg_4__0_ ( .D(n8160), .CK(GCK), .RN(n107), .Q(rd_reg[175]), 
        .QN(n809) );
  DFFRX1 rd_reg_reg_3__15_ ( .D(n1055), .CK(GCK), .RN(n109), .Q(rd_reg[206]), 
        .QN(n601) );
  DFFRX1 rd_reg_reg_3__14_ ( .D(n1039), .CK(GCK), .RN(n108), .Q(rd_reg[205]), 
        .QN(n6150) );
  DFFRX1 rd_reg_reg_3__13_ ( .D(n1023), .CK(GCK), .RN(n107), .Q(rd_reg[204]), 
        .QN(n6290) );
  DFFRX1 rd_reg_reg_3__12_ ( .D(n1007), .CK(GCK), .RN(n109), .Q(rd_reg[203]), 
        .QN(n6430) );
  DFFRX1 rd_reg_reg_3__11_ ( .D(n991), .CK(GCK), .RN(n108), .Q(rd_reg[202]), 
        .QN(n657) );
  DFFRX1 rd_reg_reg_3__10_ ( .D(n975), .CK(GCK), .RN(n107), .Q(rd_reg[201]), 
        .QN(n6710) );
  DFFRX1 rd_reg_reg_3__9_ ( .D(n959), .CK(GCK), .RN(n109), .Q(rd_reg[200]), 
        .QN(n6850) );
  DFFRX1 rd_reg_reg_3__8_ ( .D(n943), .CK(GCK), .RN(n108), .Q(rd_reg[199]), 
        .QN(n699) );
  DFFRX1 rd_reg_reg_3__2_ ( .D(n847), .CK(GCK), .RN(n107), .Q(rd_reg[193]), 
        .QN(n7830) );
  DFFRX1 rd_reg_reg_3__1_ ( .D(n8310), .CK(GCK), .RN(n109), .Q(rd_reg[192]), 
        .QN(n797) );
  DFFRX1 rd_reg_reg_3__0_ ( .D(n8150), .CK(GCK), .RN(n108), .Q(rd_reg[191]), 
        .QN(n8100) );
  DFFRX1 rd_reg_reg_2__15_ ( .D(n1054), .CK(GCK), .RN(n107), .Q(rd_reg[222]), 
        .QN(n602) );
  DFFRX1 rd_reg_reg_2__14_ ( .D(n1038), .CK(GCK), .RN(n109), .Q(rd_reg[221]), 
        .QN(n6160) );
  DFFRX1 rd_reg_reg_2__13_ ( .D(n1022), .CK(GCK), .RN(n108), .Q(rd_reg[220]), 
        .QN(n6300) );
  DFFRX1 rd_reg_reg_2__12_ ( .D(n1006), .CK(GCK), .RN(n107), .Q(rd_reg[219]), 
        .QN(n644) );
  DFFRX1 rd_reg_reg_2__11_ ( .D(n990), .CK(GCK), .RN(n109), .Q(rd_reg[218]), 
        .QN(n658) );
  DFFRX1 rd_reg_reg_2__10_ ( .D(n974), .CK(GCK), .RN(n108), .Q(rd_reg[217]), 
        .QN(n6720) );
  DFFRX1 rd_reg_reg_2__9_ ( .D(n958), .CK(GCK), .RN(n107), .Q(rd_reg[216]), 
        .QN(n6860) );
  DFFRX1 rd_reg_reg_2__8_ ( .D(n942), .CK(GCK), .RN(n109), .Q(rd_reg[215]), 
        .QN(n700) );
  DFFRX1 rd_reg_reg_2__2_ ( .D(n846), .CK(GCK), .RN(n108), .Q(rd_reg[209]), 
        .QN(n7840) );
  DFFRX1 rd_reg_reg_2__1_ ( .D(n8300), .CK(GCK), .RN(n107), .Q(rd_reg[208]), 
        .QN(n798) );
  DFFRX1 rd_reg_reg_1__15_ ( .D(n1053), .CK(GCK), .RN(n109), .Q(rd_reg[238]), 
        .QN(n603) );
  DFFRX1 rd_reg_reg_1__14_ ( .D(n1037), .CK(GCK), .RN(n108), .Q(rd_reg[237]), 
        .QN(n6170) );
  DFFRX1 rd_reg_reg_1__13_ ( .D(n1021), .CK(GCK), .RN(n107), .Q(rd_reg[236]), 
        .QN(n6310) );
  DFFRX1 rd_reg_reg_1__12_ ( .D(n1005), .CK(GCK), .RN(n109), .Q(rd_reg[235]), 
        .QN(n645) );
  DFFRX1 rd_reg_reg_1__11_ ( .D(n989), .CK(GCK), .RN(n108), .Q(rd_reg[234]), 
        .QN(n659) );
  DFFRX1 rd_reg_reg_1__10_ ( .D(n973), .CK(GCK), .RN(n107), .Q(rd_reg[233]), 
        .QN(n6730) );
  DFFRX1 rd_reg_reg_1__9_ ( .D(n957), .CK(GCK), .RN(n109), .Q(rd_reg[232]), 
        .QN(n6870) );
  DFFRX1 rd_reg_reg_1__2_ ( .D(n845), .CK(GCK), .RN(n108), .Q(rd_reg[225]), 
        .QN(n7850) );
  DFFRX1 rd_reg_reg_1__1_ ( .D(n8290), .CK(GCK), .RN(n107), .Q(rd_reg[224]), 
        .QN(n799) );
  DFFRX1 rd_reg_reg_14__4_ ( .D(n8900), .CK(GCK), .RN(n109), .Q(rd_reg[19]), 
        .QN(n744) );
  DFFRX1 rd_reg_reg_14__3_ ( .D(n8740), .CK(GCK), .RN(n108), .Q(rd_reg[18]), 
        .QN(n758) );
  DFFRX1 rd_reg_reg_14__2_ ( .D(n858), .CK(GCK), .RN(n107), .Q(rd_reg[17]), 
        .QN(n7720) );
  DFFRX1 rd_reg_reg_13__4_ ( .D(n8890), .CK(GCK), .RN(n109), .Q(rd_reg[35]), 
        .QN(n745) );
  DFFRX1 rd_reg_reg_13__3_ ( .D(n8730), .CK(GCK), .RN(n108), .Q(rd_reg[34]), 
        .QN(n759) );
  DFFRX1 rd_reg_reg_13__2_ ( .D(n857), .CK(GCK), .RN(n107), .Q(rd_reg[33]), 
        .QN(n7730) );
  DFFRX1 rd_reg_reg_12__4_ ( .D(n8880), .CK(GCK), .RN(n109), .Q(rd_reg[51]), 
        .QN(n746) );
  DFFRX1 rd_reg_reg_12__3_ ( .D(n8720), .CK(GCK), .RN(n108), .Q(rd_reg[50]), 
        .QN(n7600) );
  DFFRX1 rd_reg_reg_12__2_ ( .D(n856), .CK(GCK), .RN(n107), .Q(rd_reg[49]), 
        .QN(n7740) );
  DFFRX1 rd_reg_reg_11__4_ ( .D(n8870), .CK(GCK), .RN(n109), .Q(rd_reg[67]), 
        .QN(n747) );
  DFFRX1 rd_reg_reg_11__3_ ( .D(n8710), .CK(GCK), .RN(n108), .Q(rd_reg[66]), 
        .QN(n7610) );
  DFFRX1 rd_reg_reg_11__2_ ( .D(n855), .CK(GCK), .RN(n107), .Q(rd_reg[65]), 
        .QN(n7750) );
  DFFRX1 rd_reg_reg_10__5_ ( .D(n902), .CK(GCK), .RN(n109), .Q(rd_reg[84]), 
        .QN(n7340) );
  DFFRX1 rd_reg_reg_10__4_ ( .D(n8860), .CK(GCK), .RN(n108), .Q(rd_reg[83]), 
        .QN(n748) );
  DFFRX1 rd_reg_reg_10__3_ ( .D(n8700), .CK(GCK), .RN(n107), .Q(rd_reg[82]), 
        .QN(n7620) );
  DFFRX1 rd_reg_reg_10__2_ ( .D(n854), .CK(GCK), .RN(n109), .Q(rd_reg[81]), 
        .QN(n7760) );
  DFFRX1 rd_reg_reg_9__5_ ( .D(n901), .CK(GCK), .RN(n108), .Q(rd_reg[100]), 
        .QN(n7350) );
  DFFRX1 rd_reg_reg_9__4_ ( .D(n8850), .CK(GCK), .RN(n107), .Q(rd_reg[99]), 
        .QN(n749) );
  DFFRX1 rd_reg_reg_9__3_ ( .D(n8690), .CK(GCK), .RN(n109), .Q(rd_reg[98]), 
        .QN(n7630) );
  DFFRX1 rd_reg_reg_9__2_ ( .D(n853), .CK(GCK), .RN(n108), .Q(rd_reg[97]), 
        .QN(n7770) );
  DFFRX1 rd_reg_reg_8__5_ ( .D(n900), .CK(GCK), .RN(n107), .Q(rd_reg[116]), 
        .QN(n7360) );
  DFFRX1 rd_reg_reg_8__4_ ( .D(n8840), .CK(GCK), .RN(n109), .Q(rd_reg[115]), 
        .QN(n750) );
  DFFRX1 rd_reg_reg_8__3_ ( .D(n8680), .CK(GCK), .RN(n108), .Q(rd_reg[114]), 
        .QN(n7640) );
  DFFRX1 rd_reg_reg_8__2_ ( .D(n852), .CK(GCK), .RN(n107), .Q(rd_reg[113]), 
        .QN(n7780) );
  DFFRX1 rd_reg_reg_7__6_ ( .D(n915), .CK(GCK), .RN(n109), .Q(rd_reg[133]), 
        .QN(n7230) );
  DFFRX1 rd_reg_reg_7__5_ ( .D(n899), .CK(GCK), .RN(n108), .Q(rd_reg[132]), 
        .QN(n7370) );
  DFFRX1 rd_reg_reg_7__4_ ( .D(n8830), .CK(GCK), .RN(n107), .Q(rd_reg[131]), 
        .QN(n751) );
  DFFRX1 rd_reg_reg_7__3_ ( .D(n8670), .CK(GCK), .RN(n109), .Q(rd_reg[130]), 
        .QN(n7650) );
  DFFRX1 rd_reg_reg_7__2_ ( .D(n851), .CK(GCK), .RN(n108), .Q(rd_reg[129]), 
        .QN(n7790) );
  DFFRX1 rd_reg_reg_6__5_ ( .D(n898), .CK(GCK), .RN(n107), .Q(rd_reg[148]), 
        .QN(n7380) );
  DFFRX1 rd_reg_reg_6__4_ ( .D(n8820), .CK(GCK), .RN(n109), .Q(rd_reg[147]), 
        .QN(n752) );
  DFFRX1 rd_reg_reg_6__3_ ( .D(n8660), .CK(GCK), .RN(n108), .Q(rd_reg[146]), 
        .QN(n7660) );
  DFFRX1 rd_reg_reg_6__2_ ( .D(n850), .CK(GCK), .RN(n107), .Q(rd_reg[145]), 
        .QN(n7800) );
  DFFRX1 rd_reg_reg_5__5_ ( .D(n897), .CK(GCK), .RN(n109), .Q(rd_reg[164]), 
        .QN(n7390) );
  DFFRX1 rd_reg_reg_5__4_ ( .D(n8810), .CK(GCK), .RN(n108), .Q(rd_reg[163]), 
        .QN(n753) );
  DFFRX1 rd_reg_reg_5__3_ ( .D(n8650), .CK(GCK), .RN(n107), .Q(rd_reg[162]), 
        .QN(n7670) );
  DFFRX1 rd_reg_reg_5__2_ ( .D(n849), .CK(GCK), .RN(n109), .Q(rd_reg[161]), 
        .QN(n7810) );
  DFFRX1 rd_reg_reg_4__7_ ( .D(n928), .CK(GCK), .RN(n108), .Q(rd_reg[182]), 
        .QN(n7120) );
  DFFRX1 rd_reg_reg_4__5_ ( .D(n896), .CK(GCK), .RN(n107), .Q(rd_reg[180]), 
        .QN(n7400) );
  DFFRX1 rd_reg_reg_4__4_ ( .D(n8800), .CK(GCK), .RN(n109), .Q(rd_reg[179]), 
        .QN(n754) );
  DFFRX1 rd_reg_reg_4__3_ ( .D(n8640), .CK(GCK), .RN(n108), .Q(rd_reg[178]), 
        .QN(n7680) );
  DFFRX1 rd_reg_reg_4__2_ ( .D(n848), .CK(GCK), .RN(n107), .Q(rd_reg[177]), 
        .QN(n7820) );
  DFFRX1 rd_reg_reg_4__1_ ( .D(n8320), .CK(GCK), .RN(n109), .Q(rd_reg[176]), 
        .QN(n796) );
  DFFRX1 rd_reg_reg_3__5_ ( .D(n895), .CK(GCK), .RN(n108), .Q(rd_reg[196]), 
        .QN(n7410) );
  DFFRX1 rd_reg_reg_3__4_ ( .D(n8790), .CK(GCK), .RN(n107), .Q(rd_reg[195]), 
        .QN(n755) );
  DFFRX1 rd_reg_reg_3__3_ ( .D(n8630), .CK(GCK), .RN(n109), .Q(rd_reg[194]), 
        .QN(n7690) );
  DFFRX1 rd_reg_reg_2__5_ ( .D(n894), .CK(GCK), .RN(n108), .Q(rd_reg[212]), 
        .QN(n7420) );
  DFFRX1 rd_reg_reg_2__4_ ( .D(n8780), .CK(GCK), .RN(n107), .Q(rd_reg[211]), 
        .QN(n756) );
  DFFRX1 rd_reg_reg_2__3_ ( .D(n8620), .CK(GCK), .RN(n109), .Q(rd_reg[210]), 
        .QN(n7700) );
  DFFRX1 rd_reg_reg_1__5_ ( .D(n8930), .CK(GCK), .RN(n108), .Q(rd_reg[228]), 
        .QN(n7430) );
  DFFRX1 rd_reg_reg_1__4_ ( .D(n8770), .CK(GCK), .RN(n107), .Q(rd_reg[227]), 
        .QN(n757) );
  DFFRX1 rd_reg_reg_1__3_ ( .D(n8610), .CK(GCK), .RN(n109), .Q(rd_reg[226]), 
        .QN(n7710) );
  DFFRX1 rd_reg_reg_13__15_ ( .D(n1065), .CK(GCK), .RN(n108), .Q(rd_reg[46]), 
        .QN(n5910) );
  DFFRX1 rd_reg_reg_11__7_ ( .D(n935), .CK(GCK), .RN(n107), .Q(rd_reg[70]), 
        .QN(n705) );
  DFFRX1 rd_reg_reg_10__7_ ( .D(n934), .CK(GCK), .RN(n109), .Q(rd_reg[86]), 
        .QN(n706) );
  DFFRX1 rd_reg_reg_9__7_ ( .D(n933), .CK(GCK), .RN(n108), .Q(rd_reg[102]), 
        .QN(n707) );
  DFFRX1 rd_reg_reg_8__7_ ( .D(n932), .CK(GCK), .RN(n107), .Q(rd_reg[118]), 
        .QN(n708) );
  DFFRX1 rd_reg_reg_7__7_ ( .D(n931), .CK(GCK), .RN(n109), .Q(rd_reg[134]), 
        .QN(n709) );
  DFFRX1 rd_reg_reg_6__7_ ( .D(n930), .CK(GCK), .RN(n108), .Q(rd_reg[150]), 
        .QN(n7100) );
  DFFRX1 rd_reg_reg_1__8_ ( .D(n941), .CK(GCK), .RN(n107), .Q(rd_reg[231]), 
        .QN(n701) );
  DFFRX1 rd_reg_reg_14__15_ ( .D(n1066), .CK(GCK), .RN(n109), .Q(rd_reg[30]), 
        .QN(n5900) );
  DFFRX1 rd_reg_reg_12__15_ ( .D(n1064), .CK(GCK), .RN(n108), .Q(rd_reg[62]), 
        .QN(n5920) );
  DFFRX1 rd_reg_reg_11__15_ ( .D(n1063), .CK(GCK), .RN(n107), .Q(rd_reg[78]), 
        .QN(n5930) );
  DFFRX1 rd_reg_reg_10__15_ ( .D(n1062), .CK(GCK), .RN(n109), .Q(rd_reg[94]), 
        .QN(n594) );
  DFFRX1 rd_reg_reg_9__15_ ( .D(n1061), .CK(GCK), .RN(n108), .Q(rd_reg[110]), 
        .QN(n595) );
  DFFRX1 rd_reg_reg_8__15_ ( .D(n1060), .CK(GCK), .RN(n107), .Q(rd_reg[126]), 
        .QN(n596) );
  DFFRX1 rd_reg_reg_7__15_ ( .D(n1059), .CK(GCK), .RN(n109), .Q(rd_reg[142]), 
        .QN(n597) );
  DFFRX1 rd_reg_reg_6__15_ ( .D(n1058), .CK(GCK), .RN(n108), .Q(rd_reg[158]), 
        .QN(n598) );
  DFFRX1 rd_reg_reg_5__15_ ( .D(n1057), .CK(GCK), .RN(n107), .Q(rd_reg[174]), 
        .QN(n599) );
  DFFRX1 rd_reg_reg_4__15_ ( .D(n1056), .CK(GCK), .RN(n109), .Q(rd_reg[190]), 
        .QN(n600) );
  DFFRX1 rd_reg_reg_2__0_ ( .D(n8140), .CK(GCK), .RN(n108), .Q(rd_reg[207]), 
        .QN(n8110) );
  DFFRX1 rd_reg_reg_1__0_ ( .D(n8130), .CK(GCK), .RN(n107), .Q(rd_reg[223]), 
        .QN(n8270) );
  DFFRX1 rd_reg_reg_14__0_ ( .D(n8260), .CK(GCK), .RN(n109), .Q(rd_reg[15]) );
  DFFRX1 rd_reg_reg_13__0_ ( .D(n8250), .CK(GCK), .RN(n108), .Q(rd_reg[31]), 
        .QN(n800) );
  DFFRX1 cnt_reg_3_ ( .D(N42), .CK(GCK), .RN(n107), .Q(cnt[3]) );
  DFFRX1 cnt_reg_4_ ( .D(N43), .CK(GCK), .RN(n109), .Q(cnt[4]) );
  DFFRX1 out_buffer_reg_4__10_ ( .D(N337), .CK(GCK), .RN(n108), .Q(
        out_buffer[186]) );
  DFFRX1 out_buffer_reg_4__9_ ( .D(N336), .CK(GCK), .RN(n107), .Q(
        out_buffer[185]) );
  DFFRX1 out_buffer_reg_4__5_ ( .D(N332), .CK(GCK), .RN(n109), .Q(
        out_buffer[181]) );
  DFFRX1 out_buffer_reg_4__4_ ( .D(N331), .CK(GCK), .RN(n108), .Q(
        out_buffer[180]) );
  DFFRX1 out_buffer_reg_1__4_ ( .D(N181), .CK(GCK), .RN(n107), .Q(
        out_buffer[228]) );
  DFFRX1 out_buffer_reg_0__0_ ( .D(N127), .CK(GCK), .RN(n109), .Q(
        out_buffer[240]) );
  DFFRX1 out_buffer_reg_4__0_ ( .D(N327), .CK(GCK), .RN(n108), .Q(
        out_buffer[176]) );
  DFFRX1 out_buffer_reg_15__4_ ( .D(N881), .CK(GCK), .RN(n109), .Q(
        out_buffer[4]) );
  DFFRX1 out_buffer_reg_15__3_ ( .D(N880), .CK(GCK), .RN(n108), .Q(
        out_buffer[3]) );
  DFFRX4 r_push_reg_reg ( .D(n346), .CK(GCK), .RN(n107), .Q(r_push_reg), .QN(
        n507) );
  DFFRX1 out_buffer_reg_12__0_ ( .D(N727), .CK(GCK), .RN(n405), .Q(
        out_buffer[48]) );
  DFFRX2 out_buffer_reg_9__0_ ( .D(N577), .CK(GCK), .RN(n409), .Q(
        out_buffer[96]) );
  DFFRX1 out_buffer_reg_9__5_ ( .D(N582), .CK(GCK), .RN(n4100), .Q(
        out_buffer[101]) );
  DFFRX1 out_buffer_reg_9__8_ ( .D(N585), .CK(GCK), .RN(n4100), .Q(
        out_buffer[104]) );
  DFFRX2 out_buffer_reg_9__1_ ( .D(N578), .CK(GCK), .RN(n409), .Q(
        out_buffer[97]) );
  DFFRX1 out_buffer_reg_10__0_ ( .D(N627), .CK(GCK), .RN(n408), .Q(
        out_buffer[80]) );
  DFFRX1 out_buffer_reg_10__10_ ( .D(N637), .CK(GCK), .RN(n409), .Q(
        out_buffer[90]) );
  DFFRX1 out_buffer_reg_10__6_ ( .D(N633), .CK(GCK), .RN(n408), .Q(
        out_buffer[86]) );
  DFFRX1 out_buffer_reg_14__5_ ( .D(N832), .CK(GCK), .RN(n403), .Q(
        out_buffer[21]) );
  DFFRX1 out_buffer_reg_14__14_ ( .D(N841), .CK(GCK), .RN(n403), .Q(
        out_buffer[30]) );
  DFFRX1 out_buffer_reg_15__2_ ( .D(N879), .CK(GCK), .RN(n401), .Q(
        out_buffer[2]) );
  DFFRX1 out_buffer_reg_15__8_ ( .D(N885), .CK(GCK), .RN(n401), .Q(
        out_buffer[8]) );
  DFFRX1 out_buffer_reg_13__2_ ( .D(N779), .CK(GCK), .RN(n404), .Q(
        out_buffer[34]) );
  DFFRX1 out_buffer_reg_13__8_ ( .D(N785), .CK(GCK), .RN(n404), .Q(
        out_buffer[40]) );
  DFFRX1 out_buffer_reg_11__2_ ( .D(N679), .CK(GCK), .RN(n407), .Q(
        out_buffer[66]) );
  DFFRX1 out_buffer_reg_11__8_ ( .D(N685), .CK(GCK), .RN(n407), .Q(
        out_buffer[72]) );
  DFFRX1 out_buffer_reg_8__2_ ( .D(N529), .CK(GCK), .RN(n4110), .Q(
        out_buffer[114]) );
  DFFRX1 out_buffer_reg_8__8_ ( .D(N535), .CK(GCK), .RN(n4110), .Q(
        out_buffer[120]) );
  DFFRX1 out_buffer_reg_7__2_ ( .D(N479), .CK(GCK), .RN(n4120), .Q(
        out_buffer[130]) );
  DFFRX1 out_buffer_reg_7__8_ ( .D(N485), .CK(GCK), .RN(n4130), .Q(
        out_buffer[136]) );
  DFFRX1 out_buffer_reg_4__2_ ( .D(N329), .CK(GCK), .RN(n4170), .Q(
        out_buffer[178]) );
  DFFRX1 out_buffer_reg_4__8_ ( .D(N335), .CK(GCK), .RN(n4170), .Q(
        out_buffer[184]) );
  DFFRX1 out_buffer_reg_3__2_ ( .D(N279), .CK(GCK), .RN(n4180), .Q(
        out_buffer[194]) );
  DFFRX1 out_buffer_reg_3__8_ ( .D(N285), .CK(GCK), .RN(n4180), .Q(
        out_buffer[200]) );
  DFFRX1 out_buffer_reg_2__2_ ( .D(N229), .CK(GCK), .RN(n4190), .Q(
        out_buffer[210]) );
  DFFRX1 out_buffer_reg_2__8_ ( .D(N235), .CK(GCK), .RN(n4200), .Q(
        out_buffer[216]) );
  DFFRX1 out_buffer_reg_1__2_ ( .D(N179), .CK(GCK), .RN(n4210), .Q(
        out_buffer[226]) );
  DFFRX1 out_buffer_reg_1__8_ ( .D(N185), .CK(GCK), .RN(n4210), .Q(
        out_buffer[232]) );
  DFFRX1 out_buffer_reg_0__2_ ( .D(N129), .CK(GCK), .RN(n4220), .Q(
        out_buffer[242]) );
  DFFRX1 out_buffer_reg_0__8_ ( .D(N135), .CK(GCK), .RN(n4230), .Q(
        out_buffer[248]) );
  DFFRX1 out_buffer_reg_9__2_ ( .D(N579), .CK(GCK), .RN(n409), .Q(
        out_buffer[98]) );
  DFFRX1 out_buffer_reg_5__1_ ( .D(N378), .CK(GCK), .RN(n4150), .Q(
        out_buffer[161]) );
  DFFRX1 out_buffer_reg_5__14_ ( .D(N391), .CK(GCK), .RN(n4160), .Q(
        out_buffer[174]) );
  DFFRX1 out_buffer_reg_12__1_ ( .D(N728), .CK(GCK), .RN(n405), .Q(
        out_buffer[49]) );
  DFFRX1 out_buffer_reg_12__15_ ( .D(N742), .CK(GCK), .RN(n406), .Q(
        out_buffer[63]) );
  DFFRX1 out_buffer_reg_12__6_ ( .D(N733), .CK(GCK), .RN(n406), .Q(
        out_buffer[54]) );
  DFFRX1 out_buffer_reg_12__13_ ( .D(N740), .CK(GCK), .RN(n406), .Q(
        out_buffer[61]) );
  DFFRX1 out_buffer_reg_10__1_ ( .D(N628), .CK(GCK), .RN(n408), .Q(
        out_buffer[81]) );
  DFFRX1 out_buffer_reg_13__6_ ( .D(N783), .CK(GCK), .RN(n404), .Q(
        out_buffer[38]) );
  DFFRX1 out_buffer_reg_11__14_ ( .D(N691), .CK(GCK), .RN(n408), .Q(
        out_buffer[78]) );
  DFFRX1 out_buffer_reg_11__6_ ( .D(N683), .CK(GCK), .RN(n407), .Q(
        out_buffer[70]) );
  DFFRX1 out_buffer_reg_7__14_ ( .D(N491), .CK(GCK), .RN(n4130), .Q(
        out_buffer[142]) );
  DFFRX1 out_buffer_reg_7__6_ ( .D(N483), .CK(GCK), .RN(n4130), .Q(
        out_buffer[134]) );
  DFFRX1 out_buffer_reg_4__14_ ( .D(N341), .CK(GCK), .RN(n4180), .Q(
        out_buffer[190]) );
  DFFRX1 out_buffer_reg_4__6_ ( .D(N333), .CK(GCK), .RN(n4170), .Q(
        out_buffer[182]) );
  DFFRX1 out_buffer_reg_3__6_ ( .D(N283), .CK(GCK), .RN(n4180), .Q(
        out_buffer[198]) );
  DFFRX1 out_buffer_reg_2__14_ ( .D(N241), .CK(GCK), .RN(n4200), .Q(
        out_buffer[222]) );
  DFFRX1 out_buffer_reg_2__6_ ( .D(N233), .CK(GCK), .RN(n4200), .Q(
        out_buffer[214]) );
  DFFRX1 out_buffer_reg_1__14_ ( .D(N191), .CK(GCK), .RN(n4220), .Q(
        out_buffer[238]) );
  DFFRX1 out_buffer_reg_1__6_ ( .D(N183), .CK(GCK), .RN(n4210), .Q(
        out_buffer[230]) );
  DFFRX1 out_buffer_reg_15__12_ ( .D(N889), .CK(GCK), .RN(n402), .Q(
        out_buffer[12]) );
  DFFRX1 out_buffer_reg_15__6_ ( .D(N883), .CK(GCK), .RN(n401), .Q(
        out_buffer[6]) );
  DFFRX1 out_buffer_reg_8__15_ ( .D(N542), .CK(GCK), .RN(n4120), .Q(
        out_buffer[127]) );
  DFFRX1 out_buffer_reg_8__12_ ( .D(N539), .CK(GCK), .RN(n4120), .Q(
        out_buffer[124]) );
  DFFRX1 out_buffer_reg_8__6_ ( .D(N533), .CK(GCK), .RN(n4110), .Q(
        out_buffer[118]) );
  DFFRX1 out_buffer_reg_0__15_ ( .D(N142), .CK(GCK), .RN(n4230), .Q(
        out_buffer[255]) );
  DFFRX1 out_buffer_reg_0__12_ ( .D(N139), .CK(GCK), .RN(n4230), .Q(
        out_buffer[252]) );
  DFFRX1 out_buffer_reg_0__6_ ( .D(N133), .CK(GCK), .RN(n4230), .Q(
        out_buffer[246]) );
  DFFRX1 out_buffer_reg_5__0_ ( .D(N377), .CK(GCK), .RN(n4150), .Q(
        out_buffer[160]) );
  DFFRX1 out_buffer_reg_12__2_ ( .D(N729), .CK(GCK), .RN(n405), .Q(
        out_buffer[50]) );
  DFFRX1 out_buffer_reg_12__10_ ( .D(N737), .CK(GCK), .RN(n406), .Q(
        out_buffer[58]) );
  DFFRX1 out_buffer_reg_6__0_ ( .D(N427), .CK(GCK), .RN(n4140), .Q(
        out_buffer[144]) );
  DFFRX1 out_buffer_reg_6__1_ ( .D(N428), .CK(GCK), .RN(n4140), .Q(
        out_buffer[145]) );
  DFFRX1 out_buffer_reg_11__1_ ( .D(N678), .CK(GCK), .RN(n407), .Q(
        out_buffer[65]) );
  DFFRX1 out_buffer_reg_4__1_ ( .D(N328), .CK(GCK), .RN(n4160), .Q(
        out_buffer[177]) );
  DFFRX1 out_buffer_reg_1__1_ ( .D(N178), .CK(GCK), .RN(n4210), .Q(
        out_buffer[225]) );
  DFFRX1 out_buffer_reg_13__1_ ( .D(N778), .CK(GCK), .RN(n404), .Q(
        out_buffer[33]) );
  DFFRX1 out_buffer_reg_3__1_ ( .D(N278), .CK(GCK), .RN(n4180), .Q(
        out_buffer[193]) );
  DFFRX1 out_buffer_reg_0__1_ ( .D(N128), .CK(GCK), .RN(n4220), .Q(
        out_buffer[241]) );
  DFFRX1 out_buffer_reg_8__1_ ( .D(N528), .CK(GCK), .RN(n4110), .Q(
        out_buffer[113]) );
  DFFRX2 out_buffer_reg_14__1_ ( .D(N828), .CK(GCK), .RN(n402), .Q(
        out_buffer[17]) );
  DFFRX2 out_buffer_reg_14__0_ ( .D(N827), .CK(GCK), .RN(n402), .Q(
        out_buffer[16]) );
  DFFRX2 out_buffer_reg_15__1_ ( .D(N878), .CK(GCK), .RN(n401), .Q(
        out_buffer[1]) );
  NAND2BX2 U3 ( .AN(N226), .B(n3740), .Y(N243) );
  NAND2BX2 U4 ( .AN(N376), .B(n3750), .Y(N393) );
  OAI2BB2X1 U5 ( .B0(n3700), .B1(rd_reg[29]), .A0N(N824), .A1N(n3790), .Y(N841) );
  OAI2BB2X1 U6 ( .B0(n3660), .B1(rd_reg[254]), .A0N(N125), .A1N(n3790), .Y(
        N142) );
  OAI2BB2X1 U7 ( .B0(n355), .B1(rd_reg[126]), .A0N(N525), .A1N(n3820), .Y(N542) );
  OAI2BB2X1 U8 ( .B0(n3630), .B1(rd_reg[222]), .A0N(N225), .A1N(n3780), .Y(
        N242) );
  OAI2BB2X1 U9 ( .B0(n356), .B1(rd_reg[142]), .A0N(N475), .A1N(n3840), .Y(N492) );
  OAI2BB2X4 U10 ( .B0(n3620), .B1(rd_reg[206]), .A0N(N275), .A1N(n3770), .Y(
        N292) );
  OAI2BB2X4 U11 ( .B0(n3670), .B1(rd_reg[46]), .A0N(N775), .A1N(n3760), .Y(
        N792) );
  OAI2BB2X2 U12 ( .B0(n3730), .B1(rd_reg[94]), .A0N(N625), .A1N(n3810), .Y(
        N642) );
  OAI2BB2X2 U13 ( .B0(n3700), .B1(rd_reg[30]), .A0N(N825), .A1N(n3790), .Y(
        N842) );
  NAND2BX4 U14 ( .AN(N626), .B(n3750), .Y(N643) );
  NAND4X4 U15 ( .A(n1840), .B(data[0]), .C(data[1]), .D(data[2]), .Y(n5110) );
  NAND2BX4 U16 ( .AN(N826), .B(n3750), .Y(N843) );
  OAI2BB2X2 U17 ( .B0(n359), .B1(rd_reg[173]), .A0N(N374), .A1N(n3860), .Y(
        N391) );
  OAI2BB2X4 U18 ( .B0(n354), .B1(rd_reg[110]), .A0N(N575), .A1N(n3810), .Y(
        N592) );
  OAI2BB2X2 U19 ( .B0(n3690), .B1(rd_reg[62]), .A0N(N725), .A1N(n3860), .Y(
        N742) );
  AND2X2 U20 ( .A(data[3]), .B(n5180), .Y(n1840) );
  INVX4 U21 ( .A(n5110), .Y(n5160) );
  CLKBUFX3 U22 ( .A(n508), .Y(n504) );
  NAND2X2 U23 ( .A(n558), .B(n1900), .Y(n552) );
  XOR2X1 U24 ( .A(n5650), .B(data[13]), .Y(n5670) );
  OAI2BB2X2 U25 ( .B0(n4600), .B1(n5890), .A0N(n1830), .A1N(data[15]), .Y(
        n1067) );
  OAI2BB2XL U26 ( .B0(n3690), .B1(rd_reg[60]), .A0N(N723), .A1N(n3850), .Y(
        N740) );
  OAI2BB2XL U27 ( .B0(n359), .B1(rd_reg[172]), .A0N(N373), .A1N(n3860), .Y(
        N390) );
  OAI2BB2XL U28 ( .B0(n3640), .B1(rd_reg[238]), .A0N(N175), .A1N(n3790), .Y(
        N192) );
  OAI2BB2XL U29 ( .B0(n3600), .B1(rd_reg[190]), .A0N(N325), .A1N(n3870), .Y(
        N342) );
  OAI2BB2XL U30 ( .B0(n3710), .B1(rd_reg[78]), .A0N(N675), .A1N(n3830), .Y(
        N692) );
  OAI21X2 U31 ( .A0(n5790), .A1(n5780), .B0(n5770), .Y(n1051) );
  XNOR2X1 U32 ( .A(n5760), .B(data[15]), .Y(n5780) );
  OAI21XL U33 ( .A0(n451), .A1(n91), .B0(n79), .Y(n8750) );
  INVX3 U34 ( .A(n1930), .Y(n346) );
  AND2X2 U35 ( .A(data[4]), .B(data[5]), .Y(n89) );
  INVX3 U36 ( .A(n1019), .Y(n106) );
  INVX16 U37 ( .A(n106), .Y(n107) );
  INVX16 U38 ( .A(n106), .Y(n108) );
  INVX16 U39 ( .A(n106), .Y(n109) );
  NOR2X1 U40 ( .A(n546), .B(n559), .Y(n547) );
  AND2X6 U41 ( .A(n5160), .B(n89), .Y(n558) );
  XNOR2X1 U42 ( .A(n552), .B(data[8]), .Y(n5360) );
  OAI21X1 U43 ( .A0(n5790), .A1(n5730), .B0(n5720), .Y(n5840) );
  NAND3BXL U44 ( .AN(n546), .B(data[8]), .C(n1900), .Y(n5410) );
  AO22X4 U45 ( .A0(n90), .A1(n5890), .B0(N875), .B1(n3750), .Y(N892) );
  NAND4BX4 U46 ( .AN(n559), .B(data[10]), .C(n558), .D(data[11]), .Y(n5750) );
  NAND2BX4 U47 ( .AN(N276), .B(n3740), .Y(N293) );
  NAND2BX4 U48 ( .AN(N776), .B(n3740), .Y(N793) );
  NOR2X1 U49 ( .A(n5640), .B(n5750), .Y(n5650) );
  AO22X4 U50 ( .A0(n1930), .A1(rd_addr[10]), .B0(N58), .B1(n345), .Y(n1081) );
  NAND2BX4 U51 ( .AN(N126), .B(n3740), .Y(N143) );
  NAND2BX4 U52 ( .AN(N526), .B(n3740), .Y(N543) );
  NAND2BX4 U53 ( .AN(N876), .B(n3740), .Y(N893) );
  OAI2BB2XL U54 ( .B0(n354), .B1(rd_reg[109]), .A0N(N574), .A1N(n3810), .Y(
        N591) );
  CLKBUFX3 U55 ( .A(n503), .Y(n4710) );
  CLKAND2X3 U56 ( .A(n4680), .B(n5850), .Y(n1920) );
  NAND2X1 U57 ( .A(mode), .B(n4680), .Y(n5790) );
  NAND2BX1 U58 ( .AN(N726), .B(n3750), .Y(N743) );
  CLKBUFX2 U59 ( .A(n508), .Y(n505) );
  NOR3X1 U60 ( .A(n5750), .B(n5800), .C(n5740), .Y(n5760) );
  AO22XL U61 ( .A0(n4710), .A1(rd_reg[31]), .B0(n4690), .B1(rd_reg[15]), .Y(
        n8250) );
  AO22XL U62 ( .A0(n4680), .A1(rd_reg[224]), .B0(n498), .B1(rd_reg[240]), .Y(
        n8280) );
  AO22XL U63 ( .A0(n4680), .A1(rd_reg[225]), .B0(n498), .B1(rd_reg[241]), .Y(
        n844) );
  AO22XL U64 ( .A0(n4680), .A1(rd_reg[233]), .B0(n4730), .B1(rd_reg[249]), .Y(
        n972) );
  AO22XL U65 ( .A0(n4680), .A1(rd_reg[234]), .B0(n4750), .B1(rd_reg[250]), .Y(
        n988) );
  AO22XL U66 ( .A0(n4680), .A1(rd_reg[235]), .B0(n4740), .B1(rd_reg[251]), .Y(
        n1004) );
  AO22XL U67 ( .A0(n4680), .A1(rd_reg[237]), .B0(n498), .B1(rd_reg[253]), .Y(
        n1036) );
  CLKBUFX3 U68 ( .A(n502), .Y(n4720) );
  CLKBUFX3 U69 ( .A(n501), .Y(n4740) );
  CLKBUFX3 U70 ( .A(n501), .Y(n4750) );
  CLKBUFX3 U71 ( .A(n502), .Y(n4730) );
  INVX1 U72 ( .A(n5750), .Y(n5810) );
  AO21XL U73 ( .A0(n5820), .A1(n5810), .B0(n1920), .Y(n1830) );
  XNOR2X1 U74 ( .A(n553), .B(data[11]), .Y(n554) );
  NAND3X4 U75 ( .A(data[4]), .B(data[5]), .C(n5160), .Y(n546) );
  XNOR2XL U76 ( .A(n5160), .B(n5150), .Y(n5170) );
  NAND2XL U77 ( .A(data[0]), .B(n5180), .Y(n5260) );
  INVXL U78 ( .A(data[2]), .Y(n5220) );
  CLKINVX1 U79 ( .A(r_push_reg), .Y(n508) );
  CLKINVX2 U80 ( .A(n1930), .Y(n345) );
  AOI22XL U81 ( .A0(rd_reg[14]), .A1(n506), .B0(n1920), .B1(data[14]), .Y(
        n5770) );
  NAND3X2 U82 ( .A(n5700), .B(n5690), .C(n5680), .Y(n5830) );
  NAND2XL U83 ( .A(n1920), .B(data[12]), .Y(n5680) );
  NAND2X2 U84 ( .A(n5670), .B(n5660), .Y(n5690) );
  NAND3X2 U85 ( .A(n5630), .B(n5620), .C(n5610), .Y(n1003) );
  NAND2XL U86 ( .A(n1920), .B(data[11]), .Y(n5630) );
  NAND2X2 U87 ( .A(n5600), .B(n5660), .Y(n5620) );
  OAI211XL U88 ( .A0(out_cs[1]), .A1(out_cs[0]), .B0(n1930), .C0(n5870), .Y(
        n2800) );
  OAI32XL U89 ( .A0(n2740), .A1(out_cs[2]), .A2(out_cs[0]), .B0(n2750), .B1(
        n86), .Y(n1094) );
  NAND2XL U90 ( .A(n1920), .B(data[0]), .Y(n5280) );
  XOR2XL U91 ( .A(n5260), .B(data[1]), .Y(n5290) );
  CLKINVX1 U92 ( .A(rst), .Y(n1019) );
  INVX3 U93 ( .A(n4750), .Y(n451) );
  INVX3 U94 ( .A(n4730), .Y(n4610) );
  INVX3 U95 ( .A(n4730), .Y(n4620) );
  INVX3 U96 ( .A(n4720), .Y(n4630) );
  INVX3 U97 ( .A(n4720), .Y(n4640) );
  INVX3 U98 ( .A(n4720), .Y(n4650) );
  INVX3 U99 ( .A(n4720), .Y(n4660) );
  INVX3 U100 ( .A(n4750), .Y(n452) );
  INVX3 U101 ( .A(n4750), .Y(n453) );
  INVX3 U102 ( .A(n4750), .Y(n454) );
  INVX3 U103 ( .A(n4740), .Y(n455) );
  INVX3 U104 ( .A(n4740), .Y(n456) );
  INVX3 U105 ( .A(n4740), .Y(n457) );
  INVX3 U106 ( .A(n4740), .Y(n458) );
  INVX3 U107 ( .A(n4730), .Y(n459) );
  INVX3 U108 ( .A(n4730), .Y(n4600) );
  CLKBUFX3 U109 ( .A(n349), .Y(n3740) );
  CLKBUFX3 U110 ( .A(n348), .Y(n3820) );
  CLKBUFX3 U111 ( .A(n348), .Y(n3810) );
  CLKBUFX3 U112 ( .A(n347), .Y(n3850) );
  CLKBUFX3 U113 ( .A(n3880), .Y(n3840) );
  CLKBUFX3 U114 ( .A(n3880), .Y(n3830) );
  CLKBUFX3 U115 ( .A(n3880), .Y(n3870) );
  CLKBUFX3 U116 ( .A(n347), .Y(n3860) );
  CLKBUFX3 U117 ( .A(n351), .Y(n3760) );
  CLKBUFX3 U118 ( .A(n347), .Y(n3770) );
  CLKBUFX3 U119 ( .A(n347), .Y(n3780) );
  CLKBUFX3 U120 ( .A(n348), .Y(n3800) );
  CLKBUFX3 U121 ( .A(n348), .Y(n3790) );
  CLKBUFX3 U122 ( .A(n349), .Y(n3750) );
  CLKBUFX3 U123 ( .A(n3910), .Y(n3650) );
  CLKBUFX3 U124 ( .A(n3910), .Y(n3660) );
  CLKBUFX3 U125 ( .A(n3920), .Y(n3640) );
  CLKBUFX3 U126 ( .A(n3920), .Y(n3630) );
  CLKBUFX3 U127 ( .A(n3930), .Y(n3610) );
  CLKBUFX3 U128 ( .A(n3930), .Y(n3620) );
  CLKBUFX3 U129 ( .A(n350), .Y(n359) );
  CLKBUFX3 U130 ( .A(n394), .Y(n357) );
  CLKBUFX3 U131 ( .A(n394), .Y(n358) );
  CLKBUFX3 U132 ( .A(n347), .Y(n356) );
  CLKBUFX3 U133 ( .A(n351), .Y(n355) );
  CLKBUFX3 U134 ( .A(n350), .Y(n3600) );
  CLKBUFX3 U135 ( .A(n347), .Y(n353) );
  CLKBUFX3 U136 ( .A(n348), .Y(n354) );
  CLKBUFX3 U137 ( .A(n3890), .Y(n3700) );
  CLKBUFX3 U138 ( .A(n3890), .Y(n3690) );
  CLKBUFX3 U139 ( .A(n3900), .Y(n3680) );
  CLKBUFX3 U140 ( .A(n3900), .Y(n3670) );
  CLKBUFX3 U141 ( .A(n3930), .Y(n3730) );
  CLKBUFX3 U142 ( .A(n394), .Y(n3720) );
  CLKBUFX3 U143 ( .A(n3920), .Y(n3710) );
  INVX3 U144 ( .A(n4710), .Y(n4670) );
  INVX3 U145 ( .A(n4710), .Y(n4680) );
  INVX3 U146 ( .A(n4710), .Y(n4690) );
  CLKBUFX3 U147 ( .A(n506), .Y(n4870) );
  CLKBUFX3 U148 ( .A(n506), .Y(n4880) );
  CLKBUFX3 U149 ( .A(n506), .Y(n4890) );
  CLKBUFX3 U150 ( .A(n498), .Y(n4900) );
  CLKBUFX3 U151 ( .A(n506), .Y(n4910) );
  CLKBUFX3 U152 ( .A(n506), .Y(n4920) );
  CLKBUFX3 U153 ( .A(n506), .Y(n494) );
  CLKBUFX3 U154 ( .A(n506), .Y(n495) );
  CLKBUFX3 U155 ( .A(n497), .Y(n496) );
  CLKBUFX3 U156 ( .A(n500), .Y(n4760) );
  CLKBUFX3 U157 ( .A(n500), .Y(n4770) );
  CLKBUFX3 U158 ( .A(n500), .Y(n4780) );
  CLKBUFX3 U159 ( .A(n500), .Y(n4790) );
  CLKBUFX3 U160 ( .A(n500), .Y(n4800) );
  CLKBUFX3 U161 ( .A(n506), .Y(n4930) );
  CLKBUFX3 U162 ( .A(n499), .Y(n4810) );
  CLKBUFX3 U163 ( .A(n499), .Y(n4820) );
  CLKBUFX3 U164 ( .A(n499), .Y(n4830) );
  CLKBUFX3 U165 ( .A(n505), .Y(n4840) );
  CLKBUFX3 U166 ( .A(n498), .Y(n4850) );
  CLKBUFX3 U167 ( .A(n506), .Y(n4860) );
  CLKINVX1 U168 ( .A(n4710), .Y(n4700) );
  CLKBUFX3 U169 ( .A(n4240), .Y(n4220) );
  CLKBUFX3 U170 ( .A(n4250), .Y(n4210) );
  CLKBUFX3 U171 ( .A(n4250), .Y(n4200) );
  CLKBUFX3 U172 ( .A(n4260), .Y(n4190) );
  CLKBUFX3 U173 ( .A(n4260), .Y(n4180) );
  CLKBUFX3 U174 ( .A(n4270), .Y(n4170) );
  CLKBUFX3 U175 ( .A(n4270), .Y(n4160) );
  CLKBUFX3 U176 ( .A(n4280), .Y(n4150) );
  CLKBUFX3 U177 ( .A(n4280), .Y(n4140) );
  CLKBUFX3 U178 ( .A(n4290), .Y(n4130) );
  CLKBUFX3 U179 ( .A(n4290), .Y(n4120) );
  CLKBUFX3 U180 ( .A(n4300), .Y(n4110) );
  CLKBUFX3 U181 ( .A(n4300), .Y(n4100) );
  CLKBUFX3 U182 ( .A(n4310), .Y(n409) );
  CLKBUFX3 U183 ( .A(n4310), .Y(n408) );
  CLKBUFX3 U184 ( .A(n4320), .Y(n407) );
  CLKBUFX3 U185 ( .A(n4320), .Y(n406) );
  CLKBUFX3 U186 ( .A(n4330), .Y(n405) );
  CLKBUFX3 U187 ( .A(n4330), .Y(n404) );
  CLKBUFX3 U188 ( .A(n4340), .Y(n403) );
  CLKBUFX3 U189 ( .A(n4340), .Y(n402) );
  CLKBUFX3 U190 ( .A(n4350), .Y(n401) );
  CLKBUFX3 U191 ( .A(n4430), .Y(n400) );
  CLKBUFX3 U192 ( .A(n1019), .Y(n399) );
  CLKBUFX3 U193 ( .A(n4240), .Y(n4230) );
  CLKBUFX3 U194 ( .A(n504), .Y(n503) );
  CLKBUFX3 U195 ( .A(n507), .Y(n497) );
  CLKBUFX3 U196 ( .A(n507), .Y(n498) );
  CLKBUFX3 U197 ( .A(n504), .Y(n501) );
  CLKBUFX3 U198 ( .A(n504), .Y(n502) );
  CLKBUFX3 U199 ( .A(n349), .Y(n3910) );
  CLKBUFX3 U200 ( .A(n350), .Y(n3920) );
  CLKBUFX3 U201 ( .A(n350), .Y(n3930) );
  CLKBUFX3 U202 ( .A(n351), .Y(n394) );
  CLKBUFX3 U203 ( .A(n347), .Y(n3880) );
  CLKBUFX3 U204 ( .A(n349), .Y(n3890) );
  CLKBUFX3 U205 ( .A(n349), .Y(n3900) );
  CLKBUFX3 U206 ( .A(n507), .Y(n500) );
  CLKBUFX3 U207 ( .A(n505), .Y(n499) );
  CLKBUFX3 U208 ( .A(n449), .Y(n4260) );
  CLKBUFX3 U209 ( .A(n449), .Y(n4270) );
  CLKBUFX3 U210 ( .A(n449), .Y(n4280) );
  CLKBUFX3 U211 ( .A(n448), .Y(n4290) );
  CLKBUFX3 U212 ( .A(n448), .Y(n4300) );
  CLKBUFX3 U213 ( .A(n448), .Y(n4310) );
  CLKBUFX3 U214 ( .A(n447), .Y(n4320) );
  CLKBUFX3 U215 ( .A(n447), .Y(n4330) );
  CLKBUFX3 U216 ( .A(n447), .Y(n4340) );
  CLKBUFX3 U217 ( .A(n446), .Y(n4350) );
  CLKBUFX3 U218 ( .A(n446), .Y(n4360) );
  CLKBUFX3 U219 ( .A(n445), .Y(n4370) );
  CLKBUFX3 U220 ( .A(n445), .Y(n4380) );
  CLKBUFX3 U221 ( .A(n444), .Y(n4390) );
  CLKBUFX3 U222 ( .A(n444), .Y(n4400) );
  CLKBUFX3 U223 ( .A(n444), .Y(n4410) );
  CLKBUFX3 U224 ( .A(n4430), .Y(n4420) );
  CLKBUFX3 U225 ( .A(n450), .Y(n4240) );
  CLKBUFX3 U226 ( .A(n450), .Y(n4250) );
  XNOR2X1 U227 ( .A(n5810), .B(n5640), .Y(n5600) );
  NAND2X1 U228 ( .A(n1910), .B(n1900), .Y(n559) );
  NOR2X1 U229 ( .A(n5150), .B(n5110), .Y(n5120) );
  NOR2X1 U230 ( .A(n5220), .B(n5230), .Y(n5190) );
  CLKBUFX3 U231 ( .A(n352), .Y(n350) );
  CLKBUFX3 U232 ( .A(n352), .Y(n351) );
  CLKBUFX3 U233 ( .A(n5880), .Y(n347) );
  CLKBUFX3 U234 ( .A(n352), .Y(n349) );
  CLKBUFX3 U235 ( .A(n352), .Y(n348) );
  CLKBUFX3 U236 ( .A(n507), .Y(n506) );
  CLKBUFX3 U237 ( .A(n398), .Y(n449) );
  CLKBUFX3 U238 ( .A(n397), .Y(n448) );
  CLKBUFX3 U239 ( .A(n397), .Y(n447) );
  CLKBUFX3 U240 ( .A(n396), .Y(n446) );
  CLKBUFX3 U241 ( .A(n396), .Y(n445) );
  CLKBUFX3 U242 ( .A(n395), .Y(n444) );
  CLKBUFX3 U243 ( .A(n395), .Y(n4430) );
  CLKBUFX3 U244 ( .A(n398), .Y(n450) );
  XOR2X1 U245 ( .A(n547), .B(data[10]), .Y(n548) );
  XOR2X1 U246 ( .A(n5310), .B(data[7]), .Y(n5320) );
  NOR2X1 U247 ( .A(n5300), .B(n546), .Y(n5310) );
  NAND3BX1 U248 ( .AN(n552), .B(data[10]), .C(n1910), .Y(n553) );
  XOR2X1 U249 ( .A(n5410), .B(n5400), .Y(n5420) );
  CLKINVX1 U250 ( .A(data[9]), .Y(n5400) );
  NOR3BXL U251 ( .AN(data[14]), .B(n5800), .C(n5790), .Y(n5820) );
  AND2X2 U252 ( .A(data[7]), .B(data[6]), .Y(n1900) );
  OAI21XL U253 ( .A0(n451), .A1(n93), .B0(n63), .Y(n859) );
  AOI21X1 U254 ( .A0(n5210), .A1(n5660), .B0(n5200), .Y(n63) );
  AND2XL U255 ( .A(n1920), .B(data[2]), .Y(n5200) );
  XOR2X1 U256 ( .A(n5190), .B(data[3]), .Y(n5210) );
  AOI22XL U257 ( .A0(n5170), .A1(n5660), .B0(n1920), .B1(data[3]), .Y(n79) );
  OAI21XL U258 ( .A0(n451), .A1(n94), .B0(n95), .Y(n8910) );
  AOI21X1 U259 ( .A0(n5140), .A1(n5660), .B0(n5130), .Y(n95) );
  AND2XL U260 ( .A(n1920), .B(data[4]), .Y(n5130) );
  XOR2X1 U261 ( .A(n5120), .B(data[5]), .Y(n5140) );
  OAI21XL U262 ( .A0(n451), .A1(n87), .B0(n1110), .Y(n907) );
  AOI21X1 U263 ( .A0(n5100), .A1(n5660), .B0(n509), .Y(n1110) );
  AND2XL U264 ( .A(n1920), .B(data[5]), .Y(n509) );
  XNOR2X1 U265 ( .A(n558), .B(n5300), .Y(n5100) );
  AND2X2 U266 ( .A(data[9]), .B(data[8]), .Y(n1910) );
  NAND2BX1 U267 ( .AN(n5260), .B(data[1]), .Y(n5230) );
  NAND2X1 U268 ( .A(data[13]), .B(data[12]), .Y(n5800) );
  CLKINVX1 U269 ( .A(data[14]), .Y(n5740) );
  CLKINVX1 U270 ( .A(data[4]), .Y(n5150) );
  CLKINVX1 U271 ( .A(data[6]), .Y(n5300) );
  CLKINVX1 U272 ( .A(data[12]), .Y(n5640) );
  OAI21XL U273 ( .A0(n451), .A1(n92), .B0(n47), .Y(n8430) );
  AOI21X1 U274 ( .A0(n5250), .A1(n5660), .B0(n5240), .Y(n47) );
  AND2XL U275 ( .A(n1920), .B(data[1]), .Y(n5240) );
  XOR2X1 U276 ( .A(n5230), .B(n5220), .Y(n5250) );
  OAI22XL U277 ( .A0(n1930), .A1(n2740), .B0(n2750), .B1(n88), .Y(n1092) );
  OAI22XL U278 ( .A0(n496), .A1(n709), .B0(n451), .B1(n7100), .Y(n930) );
  OAI22XL U279 ( .A0(n496), .A1(n708), .B0(n451), .B1(n709), .Y(n931) );
  OAI22XL U280 ( .A0(n497), .A1(n707), .B0(n451), .B1(n708), .Y(n932) );
  OAI22XL U281 ( .A0(n496), .A1(n706), .B0(n451), .B1(n707), .Y(n933) );
  OAI22XL U282 ( .A0(n497), .A1(n705), .B0(n451), .B1(n706), .Y(n934) );
  OAI22XL U283 ( .A0(n4810), .A1(n704), .B0(n451), .B1(n705), .Y(n935) );
  OAI22XL U284 ( .A0(n4860), .A1(n5900), .B0(n451), .B1(n5910), .Y(n1065) );
  OAI22XL U285 ( .A0(n4870), .A1(n8100), .B0(n4600), .B1(n8110), .Y(n8140) );
  OAI22XL U286 ( .A0(n4870), .A1(n809), .B0(n4610), .B1(n8100), .Y(n8150) );
  OAI22XL U287 ( .A0(n4870), .A1(n808), .B0(n4610), .B1(n809), .Y(n8160) );
  OAI22XL U288 ( .A0(n4870), .A1(n807), .B0(n4610), .B1(n808), .Y(n8170) );
  OAI22XL U289 ( .A0(n4870), .A1(n806), .B0(n4610), .B1(n807), .Y(n8180) );
  OAI22XL U290 ( .A0(n4870), .A1(n805), .B0(n4610), .B1(n806), .Y(n8190) );
  OAI22XL U291 ( .A0(n4870), .A1(n804), .B0(n4610), .B1(n805), .Y(n8200) );
  OAI22XL U292 ( .A0(n4870), .A1(n803), .B0(n4610), .B1(n804), .Y(n8210) );
  OAI22XL U293 ( .A0(n4870), .A1(n802), .B0(n4610), .B1(n803), .Y(n8220) );
  OAI22XL U294 ( .A0(n4880), .A1(n801), .B0(n4610), .B1(n802), .Y(n8230) );
  OAI22XL U295 ( .A0(n4880), .A1(n797), .B0(n4610), .B1(n798), .Y(n8300) );
  OAI22XL U296 ( .A0(n4880), .A1(n796), .B0(n4610), .B1(n797), .Y(n8310) );
  OAI22XL U297 ( .A0(n4880), .A1(n795), .B0(n4640), .B1(n796), .Y(n8320) );
  OAI22XL U298 ( .A0(n4880), .A1(n794), .B0(n4620), .B1(n795), .Y(n8330) );
  OAI22XL U299 ( .A0(n4880), .A1(n7930), .B0(n4620), .B1(n794), .Y(n8340) );
  OAI22XL U300 ( .A0(n4880), .A1(n7920), .B0(n4620), .B1(n7930), .Y(n8350) );
  OAI22XL U301 ( .A0(n4890), .A1(n7910), .B0(n4620), .B1(n7920), .Y(n8360) );
  OAI22XL U302 ( .A0(n4890), .A1(n7900), .B0(n4620), .B1(n7910), .Y(n8370) );
  OAI22XL U303 ( .A0(n4890), .A1(n7890), .B0(n4620), .B1(n7900), .Y(n8380) );
  OAI22XL U304 ( .A0(n4890), .A1(n7880), .B0(n4620), .B1(n7890), .Y(n8390) );
  OAI22XL U305 ( .A0(n4890), .A1(n7870), .B0(n4620), .B1(n7880), .Y(n8400) );
  OAI22XL U306 ( .A0(n4890), .A1(n7860), .B0(n4620), .B1(n7870), .Y(n8410) );
  OAI22XL U307 ( .A0(n4890), .A1(n92), .B0(n4620), .B1(n7860), .Y(n8420) );
  OAI22XL U308 ( .A0(n4890), .A1(n7830), .B0(n4620), .B1(n7840), .Y(n846) );
  OAI22XL U309 ( .A0(n4900), .A1(n7820), .B0(n4620), .B1(n7830), .Y(n847) );
  OAI22XL U310 ( .A0(n4900), .A1(n7810), .B0(n4630), .B1(n7820), .Y(n848) );
  OAI22XL U311 ( .A0(n4900), .A1(n7800), .B0(n4630), .B1(n7810), .Y(n849) );
  OAI22XL U312 ( .A0(n4900), .A1(n7790), .B0(n4630), .B1(n7800), .Y(n850) );
  OAI22XL U313 ( .A0(n4900), .A1(n7780), .B0(n4630), .B1(n7790), .Y(n851) );
  OAI22XL U314 ( .A0(n4900), .A1(n7770), .B0(n4630), .B1(n7780), .Y(n852) );
  OAI22XL U315 ( .A0(n4900), .A1(n7760), .B0(n4630), .B1(n7770), .Y(n853) );
  OAI22XL U316 ( .A0(n4900), .A1(n7750), .B0(n4630), .B1(n7760), .Y(n854) );
  OAI22XL U317 ( .A0(n4900), .A1(n7740), .B0(n4630), .B1(n7750), .Y(n855) );
  OAI22XL U318 ( .A0(n4910), .A1(n7730), .B0(n4630), .B1(n7740), .Y(n856) );
  OAI22XL U319 ( .A0(n4910), .A1(n7720), .B0(n4630), .B1(n7730), .Y(n857) );
  OAI22XL U320 ( .A0(n4910), .A1(n93), .B0(n4630), .B1(n7720), .Y(n858) );
  OAI22XL U321 ( .A0(n4910), .A1(n7690), .B0(n4630), .B1(n7700), .Y(n8620) );
  OAI22XL U322 ( .A0(n4910), .A1(n7680), .B0(n4640), .B1(n7690), .Y(n8630) );
  OAI22XL U323 ( .A0(n4910), .A1(n7670), .B0(n4640), .B1(n7680), .Y(n8640) );
  OAI22XL U324 ( .A0(n4910), .A1(n7660), .B0(n4640), .B1(n7670), .Y(n8650) );
  OAI22XL U325 ( .A0(n4910), .A1(n7650), .B0(n4640), .B1(n7660), .Y(n8660) );
  OAI22XL U326 ( .A0(n4920), .A1(n7640), .B0(n4640), .B1(n7650), .Y(n8670) );
  OAI22XL U327 ( .A0(n4920), .A1(n7630), .B0(n4640), .B1(n7640), .Y(n8680) );
  OAI22XL U328 ( .A0(n4920), .A1(n7620), .B0(n4640), .B1(n7630), .Y(n8690) );
  OAI22XL U329 ( .A0(n4920), .A1(n7610), .B0(n4640), .B1(n7620), .Y(n8700) );
  OAI22XL U330 ( .A0(n4920), .A1(n7600), .B0(n4640), .B1(n7610), .Y(n8710) );
  OAI22XL U331 ( .A0(n4920), .A1(n759), .B0(n4640), .B1(n7600), .Y(n8720) );
  OAI22XL U332 ( .A0(n4920), .A1(n758), .B0(n4640), .B1(n759), .Y(n8730) );
  OAI22XL U333 ( .A0(n4920), .A1(n91), .B0(n4650), .B1(n758), .Y(n8740) );
  OAI22XL U334 ( .A0(n4930), .A1(n755), .B0(n4650), .B1(n756), .Y(n8780) );
  OAI22XL U335 ( .A0(n4930), .A1(n754), .B0(n4650), .B1(n755), .Y(n8790) );
  OAI22XL U336 ( .A0(n4930), .A1(n753), .B0(n4650), .B1(n754), .Y(n8800) );
  OAI22XL U337 ( .A0(n4930), .A1(n752), .B0(n4650), .B1(n753), .Y(n8810) );
  OAI22XL U338 ( .A0(n4930), .A1(n751), .B0(n4640), .B1(n752), .Y(n8820) );
  OAI22XL U339 ( .A0(n4930), .A1(n750), .B0(n4650), .B1(n751), .Y(n8830) );
  OAI22XL U340 ( .A0(n494), .A1(n749), .B0(n4650), .B1(n750), .Y(n8840) );
  OAI22XL U341 ( .A0(n494), .A1(n748), .B0(n4650), .B1(n749), .Y(n8850) );
  OAI22XL U342 ( .A0(n494), .A1(n747), .B0(n4650), .B1(n748), .Y(n8860) );
  OAI22XL U343 ( .A0(n494), .A1(n746), .B0(n4650), .B1(n747), .Y(n8870) );
  OAI22XL U344 ( .A0(n4930), .A1(n745), .B0(n4660), .B1(n746), .Y(n8880) );
  OAI22XL U345 ( .A0(n494), .A1(n744), .B0(n4660), .B1(n745), .Y(n8890) );
  OAI22XL U346 ( .A0(n494), .A1(n94), .B0(n4660), .B1(n744), .Y(n8900) );
  OAI22XL U347 ( .A0(n494), .A1(n7410), .B0(n4660), .B1(n7420), .Y(n894) );
  OAI22XL U348 ( .A0(n495), .A1(n7400), .B0(n4660), .B1(n7410), .Y(n895) );
  OAI22XL U349 ( .A0(n495), .A1(n7390), .B0(n4660), .B1(n7400), .Y(n896) );
  OAI22XL U350 ( .A0(n495), .A1(n7380), .B0(n4660), .B1(n7390), .Y(n897) );
  OAI22XL U351 ( .A0(n495), .A1(n7370), .B0(n4650), .B1(n7380), .Y(n898) );
  OAI22XL U352 ( .A0(n497), .A1(n7360), .B0(n4660), .B1(n7370), .Y(n899) );
  OAI22XL U353 ( .A0(n495), .A1(n7350), .B0(n4660), .B1(n7360), .Y(n900) );
  OAI22XL U354 ( .A0(n494), .A1(n7340), .B0(n4650), .B1(n7350), .Y(n901) );
  OAI22XL U355 ( .A0(n4930), .A1(n7330), .B0(n4660), .B1(n7340), .Y(n902) );
  OAI22XL U356 ( .A0(n495), .A1(n7220), .B0(n4660), .B1(n7230), .Y(n915) );
  OAI22XL U357 ( .A0(n496), .A1(n7110), .B0(n4660), .B1(n7120), .Y(n928) );
  OAI22XL U358 ( .A0(n497), .A1(n7100), .B0(n455), .B1(n7110), .Y(n929) );
  OAI22XL U359 ( .A0(n4840), .A1(n703), .B0(n452), .B1(n704), .Y(n936) );
  OAI22XL U360 ( .A0(n4840), .A1(n702), .B0(n452), .B1(n703), .Y(n937) );
  OAI22XL U361 ( .A0(n4840), .A1(n699), .B0(n452), .B1(n700), .Y(n942) );
  OAI22XL U362 ( .A0(n4840), .A1(n698), .B0(n452), .B1(n699), .Y(n943) );
  OAI22XL U363 ( .A0(n4840), .A1(n697), .B0(n452), .B1(n698), .Y(n944) );
  OAI22XL U364 ( .A0(n4760), .A1(n696), .B0(n452), .B1(n697), .Y(n945) );
  OAI22XL U365 ( .A0(n4760), .A1(n695), .B0(n452), .B1(n696), .Y(n946) );
  OAI22XL U366 ( .A0(n4760), .A1(n694), .B0(n452), .B1(n695), .Y(n947) );
  OAI22XL U367 ( .A0(n4760), .A1(n6930), .B0(n452), .B1(n694), .Y(n948) );
  OAI22XL U368 ( .A0(n4760), .A1(n6920), .B0(n453), .B1(n6930), .Y(n949) );
  OAI22XL U369 ( .A0(n4760), .A1(n6910), .B0(n452), .B1(n6920), .Y(n950) );
  OAI22XL U370 ( .A0(n4760), .A1(n6900), .B0(n453), .B1(n6910), .Y(n951) );
  OAI22XL U371 ( .A0(n4760), .A1(n6890), .B0(n452), .B1(n6900), .Y(n952) );
  OAI22XL U372 ( .A0(n4760), .A1(n6880), .B0(n453), .B1(n6890), .Y(n953) );
  OAI22XL U373 ( .A0(n4770), .A1(n6850), .B0(n453), .B1(n6860), .Y(n958) );
  OAI22XL U374 ( .A0(n4770), .A1(n6840), .B0(n453), .B1(n6850), .Y(n959) );
  OAI22XL U375 ( .A0(n4770), .A1(n6830), .B0(n453), .B1(n6840), .Y(n960) );
  OAI22XL U376 ( .A0(n4770), .A1(n6820), .B0(n453), .B1(n6830), .Y(n961) );
  OAI22XL U377 ( .A0(n4770), .A1(n6810), .B0(n453), .B1(n6820), .Y(n962) );
  OAI22XL U378 ( .A0(n4770), .A1(n6800), .B0(n453), .B1(n6810), .Y(n963) );
  OAI22XL U379 ( .A0(n4770), .A1(n6790), .B0(n453), .B1(n6800), .Y(n964) );
  OAI22XL U380 ( .A0(n4780), .A1(n6780), .B0(n453), .B1(n6790), .Y(n965) );
  OAI22XL U381 ( .A0(n4780), .A1(n6770), .B0(n453), .B1(n6780), .Y(n966) );
  OAI22XL U382 ( .A0(n4780), .A1(n6760), .B0(n454), .B1(n6770), .Y(n967) );
  OAI22XL U383 ( .A0(n4780), .A1(n6750), .B0(n454), .B1(n6760), .Y(n968) );
  OAI22XL U384 ( .A0(n4780), .A1(n6740), .B0(n454), .B1(n6750), .Y(n969) );
  OAI22XL U385 ( .A0(n4780), .A1(n6710), .B0(n454), .B1(n6720), .Y(n974) );
  OAI22XL U386 ( .A0(n4780), .A1(n6700), .B0(n454), .B1(n6710), .Y(n975) );
  OAI22XL U387 ( .A0(n4790), .A1(n6690), .B0(n454), .B1(n6700), .Y(n976) );
  OAI22XL U388 ( .A0(n4790), .A1(n6680), .B0(n454), .B1(n6690), .Y(n977) );
  OAI22XL U389 ( .A0(n4790), .A1(n6670), .B0(n454), .B1(n6680), .Y(n978) );
  OAI22XL U390 ( .A0(n4790), .A1(n6660), .B0(n454), .B1(n6670), .Y(n979) );
  OAI22XL U391 ( .A0(n4790), .A1(n6650), .B0(n455), .B1(n6660), .Y(n980) );
  OAI22XL U392 ( .A0(n4790), .A1(n6640), .B0(n454), .B1(n6650), .Y(n981) );
  OAI22XL U393 ( .A0(n4790), .A1(n6630), .B0(n454), .B1(n6640), .Y(n982) );
  OAI22XL U394 ( .A0(n4790), .A1(n6620), .B0(n455), .B1(n6630), .Y(n983) );
  OAI22XL U395 ( .A0(n4790), .A1(n6610), .B0(n455), .B1(n6620), .Y(n984) );
  OAI22XL U396 ( .A0(n4800), .A1(n6600), .B0(n455), .B1(n6610), .Y(n985) );
  OAI22XL U397 ( .A0(n4800), .A1(n657), .B0(n455), .B1(n658), .Y(n990) );
  OAI22XL U398 ( .A0(n4800), .A1(n656), .B0(n455), .B1(n657), .Y(n991) );
  OAI22XL U399 ( .A0(n4800), .A1(n655), .B0(n455), .B1(n656), .Y(n992) );
  OAI22XL U400 ( .A0(n4800), .A1(n654), .B0(n455), .B1(n655), .Y(n993) );
  OAI22XL U401 ( .A0(n4800), .A1(n653), .B0(n455), .B1(n654), .Y(n994) );
  OAI22XL U402 ( .A0(n4800), .A1(n652), .B0(n455), .B1(n653), .Y(n995) );
  OAI22XL U403 ( .A0(n4810), .A1(n651), .B0(n456), .B1(n652), .Y(n996) );
  OAI22XL U404 ( .A0(n4810), .A1(n650), .B0(n456), .B1(n651), .Y(n997) );
  OAI22XL U405 ( .A0(n4810), .A1(n649), .B0(n456), .B1(n650), .Y(n998) );
  OAI22XL U406 ( .A0(n4930), .A1(n648), .B0(n456), .B1(n649), .Y(n999) );
  OAI22XL U407 ( .A0(n4810), .A1(n647), .B0(n456), .B1(n648), .Y(n1000) );
  OAI22XL U408 ( .A0(n4810), .A1(n646), .B0(n456), .B1(n647), .Y(n1001) );
  OAI22XL U409 ( .A0(n4810), .A1(n6430), .B0(n456), .B1(n644), .Y(n1006) );
  OAI22XL U410 ( .A0(n4820), .A1(n6420), .B0(n456), .B1(n6430), .Y(n1007) );
  OAI22XL U411 ( .A0(n4820), .A1(n6410), .B0(n456), .B1(n6420), .Y(n1008) );
  OAI22XL U412 ( .A0(n4820), .A1(n6400), .B0(n456), .B1(n6410), .Y(n1009) );
  OAI22XL U413 ( .A0(n4820), .A1(n6390), .B0(n456), .B1(n6400), .Y(n1010) );
  OAI22XL U414 ( .A0(n4820), .A1(n6380), .B0(n457), .B1(n6390), .Y(n1011) );
  OAI22XL U415 ( .A0(n4820), .A1(n6370), .B0(n457), .B1(n6380), .Y(n1012) );
  OAI22XL U416 ( .A0(n4820), .A1(n6360), .B0(n457), .B1(n6370), .Y(n1013) );
  OAI22XL U417 ( .A0(n4820), .A1(n6350), .B0(n457), .B1(n6360), .Y(n1014) );
  OAI22XL U418 ( .A0(n4820), .A1(n6340), .B0(n457), .B1(n6350), .Y(n1015) );
  OAI22XL U419 ( .A0(n4830), .A1(n6330), .B0(n457), .B1(n6340), .Y(n1016) );
  OAI22XL U420 ( .A0(n4830), .A1(n6320), .B0(n457), .B1(n6330), .Y(n1017) );
  OAI22XL U421 ( .A0(n4830), .A1(n6290), .B0(n457), .B1(n6300), .Y(n1022) );
  OAI22XL U422 ( .A0(n4830), .A1(n6280), .B0(n457), .B1(n6290), .Y(n1023) );
  OAI22XL U423 ( .A0(n4830), .A1(n6270), .B0(n457), .B1(n6280), .Y(n1024) );
  OAI22XL U424 ( .A0(n4830), .A1(n6260), .B0(n457), .B1(n6270), .Y(n1025) );
  OAI22XL U425 ( .A0(n4830), .A1(n6250), .B0(n458), .B1(n6260), .Y(n1026) );
  OAI22XL U426 ( .A0(n4840), .A1(n6240), .B0(n458), .B1(n6250), .Y(n1027) );
  OAI22XL U427 ( .A0(n4840), .A1(n6230), .B0(n458), .B1(n6240), .Y(n1028) );
  OAI22XL U428 ( .A0(n4840), .A1(n6220), .B0(n458), .B1(n6230), .Y(n1029) );
  OAI22XL U429 ( .A0(n4840), .A1(n6210), .B0(n458), .B1(n6220), .Y(n1030) );
  OAI22XL U430 ( .A0(n4840), .A1(n6200), .B0(n458), .B1(n6210), .Y(n1031) );
  OAI22XL U431 ( .A0(n4840), .A1(n6190), .B0(n458), .B1(n6200), .Y(n1032) );
  OAI22XL U432 ( .A0(n4840), .A1(n6180), .B0(n458), .B1(n6190), .Y(n1033) );
  OAI22XL U433 ( .A0(n497), .A1(n6150), .B0(n458), .B1(n6160), .Y(n1038) );
  OAI22XL U434 ( .A0(n507), .A1(n6140), .B0(n458), .B1(n6150), .Y(n1039) );
  OAI22XL U435 ( .A0(n507), .A1(n6130), .B0(n458), .B1(n6140), .Y(n1040) );
  OAI22XL U436 ( .A0(n507), .A1(n6120), .B0(n459), .B1(n6130), .Y(n1041) );
  OAI22XL U437 ( .A0(n507), .A1(n6110), .B0(n459), .B1(n6120), .Y(n1042) );
  OAI22XL U438 ( .A0(n507), .A1(n6100), .B0(n459), .B1(n6110), .Y(n1043) );
  OAI22XL U439 ( .A0(n507), .A1(n609), .B0(n459), .B1(n6100), .Y(n1044) );
  OAI22XL U440 ( .A0(n507), .A1(n608), .B0(n459), .B1(n609), .Y(n1045) );
  OAI22XL U441 ( .A0(n507), .A1(n607), .B0(n459), .B1(n608), .Y(n1046) );
  OAI22XL U442 ( .A0(n4850), .A1(n606), .B0(n459), .B1(n607), .Y(n1047) );
  OAI22XL U443 ( .A0(n4850), .A1(n605), .B0(n459), .B1(n606), .Y(n1048) );
  OAI22XL U444 ( .A0(n4850), .A1(n604), .B0(n459), .B1(n605), .Y(n1049) );
  OAI22XL U445 ( .A0(n4850), .A1(n601), .B0(n459), .B1(n602), .Y(n1054) );
  OAI22XL U446 ( .A0(n4850), .A1(n600), .B0(n459), .B1(n601), .Y(n1055) );
  OAI22XL U447 ( .A0(n4850), .A1(n599), .B0(n4600), .B1(n600), .Y(n1056) );
  OAI22XL U448 ( .A0(n4850), .A1(n598), .B0(n4600), .B1(n599), .Y(n1057) );
  OAI22XL U449 ( .A0(n4860), .A1(n597), .B0(n4600), .B1(n598), .Y(n1058) );
  OAI22XL U450 ( .A0(n4860), .A1(n596), .B0(n4600), .B1(n597), .Y(n1059) );
  OAI22XL U451 ( .A0(n4860), .A1(n595), .B0(n4600), .B1(n596), .Y(n1060) );
  OAI22XL U452 ( .A0(n4860), .A1(n594), .B0(n4600), .B1(n595), .Y(n1061) );
  OAI22XL U453 ( .A0(n4860), .A1(n5930), .B0(n4600), .B1(n594), .Y(n1062) );
  OAI22XL U454 ( .A0(n4860), .A1(n5920), .B0(n4600), .B1(n5930), .Y(n1063) );
  OAI22XL U455 ( .A0(n4860), .A1(n5910), .B0(n4600), .B1(n5920), .Y(n1064) );
  OAI22XL U456 ( .A0(n4840), .A1(n5890), .B0(n4600), .B1(n5900), .Y(n1066) );
  OAI22XL U457 ( .A0(n495), .A1(n7320), .B0(n4670), .B1(n7330), .Y(n903) );
  OAI22XL U458 ( .A0(n507), .A1(n7310), .B0(n4670), .B1(n7320), .Y(n904) );
  OAI22XL U459 ( .A0(n507), .A1(n7300), .B0(n4670), .B1(n7310), .Y(n905) );
  OAI22XL U460 ( .A0(n495), .A1(n87), .B0(n4670), .B1(n7300), .Y(n906) );
  OAI22XL U461 ( .A0(n496), .A1(n7270), .B0(n4670), .B1(n7280), .Y(n910) );
  OAI22XL U462 ( .A0(n496), .A1(n7260), .B0(n4670), .B1(n7270), .Y(n911) );
  OAI22XL U463 ( .A0(n496), .A1(n7240), .B0(n4670), .B1(n7250), .Y(n913) );
  OAI22XL U464 ( .A0(n494), .A1(n7230), .B0(n4670), .B1(n7240), .Y(n914) );
  OAI22XL U465 ( .A0(n507), .A1(n7200), .B0(n4670), .B1(n7210), .Y(n917) );
  OAI22XL U466 ( .A0(n497), .A1(n7170), .B0(n4670), .B1(n7180), .Y(n920) );
  OAI22XL U467 ( .A0(n507), .A1(n7130), .B0(n4670), .B1(n7140), .Y(n926) );
  OAI22XL U468 ( .A0(n506), .A1(n7250), .B0(n4680), .B1(n7260), .Y(n912) );
  OAI22XL U469 ( .A0(n496), .A1(n7210), .B0(n4680), .B1(n7220), .Y(n916) );
  OAI22XL U470 ( .A0(n496), .A1(n7190), .B0(n4680), .B1(n7200), .Y(n918) );
  OAI22XL U471 ( .A0(n506), .A1(n7180), .B0(n4680), .B1(n7190), .Y(n919) );
  OAI22XL U472 ( .A0(n506), .A1(n7160), .B0(n4680), .B1(n7170), .Y(n921) );
  OAI22XL U473 ( .A0(n497), .A1(n7120), .B0(n4680), .B1(n7130), .Y(n927) );
  INVX3 U474 ( .A(n5790), .Y(n5660) );
  CLKINVX1 U475 ( .A(n1075), .Y(n5870) );
  CLKBUFX3 U476 ( .A(n5880), .Y(n352) );
  CLKBUFX3 U477 ( .A(n107), .Y(n398) );
  CLKBUFX3 U478 ( .A(n108), .Y(n397) );
  CLKBUFX3 U479 ( .A(n109), .Y(n396) );
  CLKBUFX3 U480 ( .A(n107), .Y(n395) );
  AOI22X1 U481 ( .A0(n1920), .A1(data[13]), .B0(n497), .B1(rd_reg[13]), .Y(
        n5720) );
  XOR2X1 U482 ( .A(n5710), .B(n5740), .Y(n5730) );
  NOR2X1 U483 ( .A(n5800), .B(n5750), .Y(n5710) );
  OAI2BB2XL U484 ( .B0(n359), .B1(rd_reg[174]), .A0N(N375), .A1N(n3860), .Y(
        N392) );
  OAI2BB2XL U485 ( .B0(n358), .B1(rd_reg[158]), .A0N(N425), .A1N(n3850), .Y(
        N442) );
  NAND3X1 U486 ( .A(n557), .B(n556), .C(n555), .Y(n987) );
  NAND2BX1 U487 ( .AN(n4690), .B(rd_reg[10]), .Y(n557) );
  NAND2X1 U488 ( .A(n1920), .B(data[10]), .Y(n555) );
  NAND2X1 U489 ( .A(n554), .B(n5660), .Y(n556) );
  NAND3X1 U490 ( .A(n545), .B(n544), .C(n5430), .Y(n955) );
  NAND2BX1 U491 ( .AN(n4690), .B(rd_reg[8]), .Y(n545) );
  NAND2X1 U492 ( .A(n1920), .B(data[8]), .Y(n5430) );
  NAND2X1 U493 ( .A(n5420), .B(n5660), .Y(n544) );
  NAND2BX1 U494 ( .AN(N176), .B(n3740), .Y(N193) );
  NAND2BX1 U495 ( .AN(N326), .B(n3740), .Y(N343) );
  NAND2BX1 U496 ( .AN(N476), .B(n3740), .Y(N493) );
  NAND2BX1 U497 ( .AN(N676), .B(n3740), .Y(N693) );
  NAND2BX1 U498 ( .AN(N426), .B(n3750), .Y(N443) );
  NAND2BX1 U499 ( .AN(N576), .B(n3750), .Y(N593) );
  NAND3X1 U500 ( .A(n5390), .B(n5380), .C(n5370), .Y(n939) );
  NAND2BX1 U501 ( .AN(n4690), .B(rd_reg[7]), .Y(n5390) );
  NAND2X1 U502 ( .A(n1920), .B(data[7]), .Y(n5370) );
  NAND2X1 U503 ( .A(n5360), .B(n5660), .Y(n5380) );
  NAND3X1 U504 ( .A(n551), .B(n550), .C(n549), .Y(n971) );
  NAND2BX1 U505 ( .AN(n4700), .B(rd_reg[9]), .Y(n551) );
  NAND2X1 U506 ( .A(n1920), .B(data[9]), .Y(n549) );
  NAND2X1 U507 ( .A(n548), .B(n5660), .Y(n550) );
  NAND2BX1 U508 ( .AN(n4690), .B(rd_reg[12]), .Y(n5700) );
  NAND3X1 U509 ( .A(n5350), .B(n5340), .C(n5330), .Y(n923) );
  NAND2BX1 U510 ( .AN(n4690), .B(rd_reg[6]), .Y(n5350) );
  NAND2X1 U511 ( .A(n1920), .B(data[6]), .Y(n5330) );
  NAND2X1 U512 ( .A(n5320), .B(n5660), .Y(n5340) );
  NAND2BX1 U513 ( .AN(n4690), .B(rd_reg[11]), .Y(n5610) );
  OAI211X1 U514 ( .A0(n5790), .A1(n5290), .B0(n5280), .C0(n5270), .Y(n5860) );
  NAND2BX1 U515 ( .AN(n4690), .B(rd_reg[0]), .Y(n5270) );
  OAI2BB2XL U516 ( .B0(n3730), .B1(rd_reg[14]), .A0N(N874), .A1N(n3760), .Y(
        N891) );
  OAI2BB2XL U517 ( .B0(n3730), .B1(rd_reg[13]), .A0N(N873), .A1N(n3760), .Y(
        N890) );
  OAI2BB2XL U518 ( .B0(n3740), .B1(rd_reg[12]), .A0N(N872), .A1N(n3770), .Y(
        N889) );
  OAI2BB2XL U519 ( .B0(n3730), .B1(rd_reg[11]), .A0N(N871), .A1N(n3770), .Y(
        N888) );
  OAI2BB2XL U520 ( .B0(n3740), .B1(rd_reg[10]), .A0N(N870), .A1N(n3780), .Y(
        N887) );
  OAI2BB2XL U521 ( .B0(n3730), .B1(rd_reg[9]), .A0N(N869), .A1N(n3780), .Y(
        N886) );
  OAI2BB2XL U522 ( .B0(n3640), .B1(rd_reg[237]), .A0N(N174), .A1N(n3790), .Y(
        N191) );
  OAI2BB2XL U523 ( .B0(n3650), .B1(rd_reg[236]), .A0N(N173), .A1N(n3790), .Y(
        N190) );
  OAI2BB2XL U524 ( .B0(n3650), .B1(rd_reg[235]), .A0N(N172), .A1N(n3800), .Y(
        N189) );
  OAI2BB2XL U525 ( .B0(n3650), .B1(rd_reg[234]), .A0N(N171), .A1N(n3800), .Y(
        N188) );
  OAI2BB2XL U526 ( .B0(n3650), .B1(rd_reg[233]), .A0N(N170), .A1N(n3800), .Y(
        N187) );
  OAI2BB2XL U527 ( .B0(n3650), .B1(rd_reg[232]), .A0N(N169), .A1N(n3800), .Y(
        N186) );
  OAI2BB2XL U528 ( .B0(n3660), .B1(rd_reg[253]), .A0N(N124), .A1N(n3790), .Y(
        N141) );
  OAI2BB2XL U529 ( .B0(n3660), .B1(rd_reg[252]), .A0N(N123), .A1N(n3790), .Y(
        N140) );
  OAI2BB2XL U530 ( .B0(n3660), .B1(rd_reg[251]), .A0N(N122), .A1N(n3780), .Y(
        N139) );
  OAI2BB2XL U531 ( .B0(n3660), .B1(rd_reg[250]), .A0N(N121), .A1N(n3780), .Y(
        N138) );
  OAI2BB2XL U532 ( .B0(n3660), .B1(rd_reg[249]), .A0N(N120), .A1N(n3780), .Y(
        N137) );
  OAI2BB2XL U533 ( .B0(n3660), .B1(rd_reg[248]), .A0N(N119), .A1N(n3780), .Y(
        N136) );
  OAI2BB2XL U534 ( .B0(n3630), .B1(rd_reg[221]), .A0N(N224), .A1N(n3780), .Y(
        N241) );
  OAI2BB2XL U535 ( .B0(n3630), .B1(rd_reg[220]), .A0N(N223), .A1N(n3780), .Y(
        N240) );
  OAI2BB2XL U536 ( .B0(n3630), .B1(rd_reg[219]), .A0N(N222), .A1N(n3780), .Y(
        N239) );
  OAI2BB2XL U537 ( .B0(n3630), .B1(rd_reg[218]), .A0N(N221), .A1N(n3780), .Y(
        N238) );
  OAI2BB2XL U538 ( .B0(n3630), .B1(rd_reg[217]), .A0N(N220), .A1N(n3780), .Y(
        N237) );
  OAI2BB2XL U539 ( .B0(n3640), .B1(rd_reg[216]), .A0N(N219), .A1N(n3780), .Y(
        N236) );
  OAI2BB2XL U540 ( .B0(n3620), .B1(rd_reg[205]), .A0N(N274), .A1N(n3760), .Y(
        N291) );
  OAI2BB2XL U541 ( .B0(n3620), .B1(rd_reg[204]), .A0N(N273), .A1N(n3760), .Y(
        N290) );
  OAI2BB2XL U542 ( .B0(n3620), .B1(rd_reg[203]), .A0N(N272), .A1N(n3760), .Y(
        N289) );
  OAI2BB2XL U543 ( .B0(n3620), .B1(rd_reg[202]), .A0N(N271), .A1N(n3760), .Y(
        N288) );
  OAI2BB2XL U544 ( .B0(n3620), .B1(rd_reg[201]), .A0N(N270), .A1N(n3770), .Y(
        N287) );
  OAI2BB2XL U545 ( .B0(n3620), .B1(rd_reg[200]), .A0N(N269), .A1N(n3770), .Y(
        N286) );
  OAI2BB2XL U546 ( .B0(n3600), .B1(rd_reg[189]), .A0N(N324), .A1N(n3870), .Y(
        N341) );
  OAI2BB2XL U547 ( .B0(n3610), .B1(rd_reg[188]), .A0N(N323), .A1N(n3870), .Y(
        N340) );
  OAI2BB2XL U548 ( .B0(n3610), .B1(rd_reg[187]), .A0N(N322), .A1N(n3870), .Y(
        N339) );
  OAI2BB2XL U549 ( .B0(n3610), .B1(rd_reg[186]), .A0N(N321), .A1N(n3870), .Y(
        N338) );
  OAI2BB2XL U550 ( .B0(n3610), .B1(rd_reg[185]), .A0N(N320), .A1N(n3760), .Y(
        N337) );
  OAI2BB2XL U551 ( .B0(n3610), .B1(rd_reg[184]), .A0N(N319), .A1N(n3600), .Y(
        N336) );
  OAI2BB2XL U552 ( .B0(n359), .B1(rd_reg[171]), .A0N(N372), .A1N(n3860), .Y(
        N389) );
  OAI2BB2XL U553 ( .B0(n359), .B1(rd_reg[170]), .A0N(N371), .A1N(n3860), .Y(
        N388) );
  OAI2BB2XL U554 ( .B0(n359), .B1(rd_reg[169]), .A0N(N370), .A1N(n3860), .Y(
        N387) );
  OAI2BB2XL U555 ( .B0(n359), .B1(rd_reg[168]), .A0N(N369), .A1N(n3860), .Y(
        N386) );
  OAI2BB2XL U556 ( .B0(n358), .B1(rd_reg[157]), .A0N(N424), .A1N(n3850), .Y(
        N441) );
  OAI2BB2XL U557 ( .B0(n358), .B1(rd_reg[156]), .A0N(N423), .A1N(n3850), .Y(
        N440) );
  OAI2BB2XL U558 ( .B0(n358), .B1(rd_reg[155]), .A0N(N422), .A1N(n3850), .Y(
        N439) );
  OAI2BB2XL U559 ( .B0(n358), .B1(rd_reg[154]), .A0N(N421), .A1N(n3850), .Y(
        N438) );
  OAI2BB2XL U560 ( .B0(n358), .B1(rd_reg[153]), .A0N(N420), .A1N(n3850), .Y(
        N437) );
  OAI2BB2XL U561 ( .B0(n358), .B1(rd_reg[152]), .A0N(N419), .A1N(n3850), .Y(
        N436) );
  OAI2BB2XL U562 ( .B0(n356), .B1(rd_reg[141]), .A0N(N474), .A1N(n3840), .Y(
        N491) );
  OAI2BB2XL U563 ( .B0(n356), .B1(rd_reg[140]), .A0N(N473), .A1N(n3840), .Y(
        N490) );
  OAI2BB2XL U564 ( .B0(n357), .B1(rd_reg[139]), .A0N(N472), .A1N(n3840), .Y(
        N489) );
  OAI2BB2XL U565 ( .B0(n357), .B1(rd_reg[138]), .A0N(N471), .A1N(n3840), .Y(
        N488) );
  OAI2BB2XL U566 ( .B0(n357), .B1(rd_reg[137]), .A0N(N470), .A1N(n3840), .Y(
        N487) );
  OAI2BB2XL U567 ( .B0(n357), .B1(rd_reg[136]), .A0N(N469), .A1N(n3840), .Y(
        N486) );
  OAI2BB2XL U568 ( .B0(n355), .B1(rd_reg[125]), .A0N(N524), .A1N(n3830), .Y(
        N541) );
  OAI2BB2XL U569 ( .B0(n355), .B1(rd_reg[124]), .A0N(N523), .A1N(n3830), .Y(
        N540) );
  OAI2BB2XL U570 ( .B0(n355), .B1(rd_reg[123]), .A0N(N522), .A1N(n3830), .Y(
        N539) );
  OAI2BB2XL U571 ( .B0(n355), .B1(rd_reg[122]), .A0N(N521), .A1N(n3830), .Y(
        N538) );
  OAI2BB2XL U572 ( .B0(n355), .B1(rd_reg[121]), .A0N(N520), .A1N(n3830), .Y(
        N537) );
  OAI2BB2XL U573 ( .B0(n355), .B1(rd_reg[120]), .A0N(N519), .A1N(n3830), .Y(
        N536) );
  OAI2BB2XL U574 ( .B0(n354), .B1(rd_reg[108]), .A0N(N573), .A1N(n3810), .Y(
        N590) );
  OAI2BB2XL U575 ( .B0(n354), .B1(rd_reg[107]), .A0N(N572), .A1N(n3810), .Y(
        N589) );
  OAI2BB2XL U576 ( .B0(n354), .B1(rd_reg[106]), .A0N(N571), .A1N(n3820), .Y(
        N588) );
  OAI2BB2XL U577 ( .B0(n354), .B1(rd_reg[105]), .A0N(N570), .A1N(n3820), .Y(
        N587) );
  OAI2BB2XL U578 ( .B0(n354), .B1(rd_reg[104]), .A0N(N569), .A1N(n3820), .Y(
        N586) );
  OAI2BB2XL U579 ( .B0(n3720), .B1(rd_reg[93]), .A0N(N624), .A1N(n3810), .Y(
        N641) );
  OAI2BB2XL U580 ( .B0(n3720), .B1(rd_reg[92]), .A0N(N623), .A1N(n3800), .Y(
        N640) );
  OAI2BB2XL U581 ( .B0(n3600), .B1(rd_reg[91]), .A0N(N622), .A1N(n3770), .Y(
        N639) );
  OAI2BB2XL U582 ( .B0(n353), .B1(rd_reg[90]), .A0N(N621), .A1N(n3840), .Y(
        N638) );
  OAI2BB2XL U583 ( .B0(n353), .B1(rd_reg[89]), .A0N(N620), .A1N(n3800), .Y(
        N637) );
  OAI2BB2XL U584 ( .B0(n353), .B1(rd_reg[88]), .A0N(N619), .A1N(n3810), .Y(
        N636) );
  OAI2BB2XL U585 ( .B0(n3710), .B1(rd_reg[77]), .A0N(N674), .A1N(n3830), .Y(
        N691) );
  OAI2BB2XL U586 ( .B0(n3710), .B1(rd_reg[76]), .A0N(N673), .A1N(n3830), .Y(
        N690) );
  OAI2BB2XL U587 ( .B0(n3720), .B1(rd_reg[75]), .A0N(N672), .A1N(n3830), .Y(
        N689) );
  OAI2BB2XL U588 ( .B0(n3720), .B1(rd_reg[74]), .A0N(N671), .A1N(n3830), .Y(
        N688) );
  OAI2BB2XL U589 ( .B0(n3720), .B1(rd_reg[73]), .A0N(N670), .A1N(n3820), .Y(
        N687) );
  OAI2BB2XL U590 ( .B0(n3720), .B1(rd_reg[72]), .A0N(N669), .A1N(n3820), .Y(
        N686) );
  OAI2BB2XL U591 ( .B0(n3690), .B1(rd_reg[61]), .A0N(N724), .A1N(n3860), .Y(
        N741) );
  OAI2BB2XL U592 ( .B0(n3690), .B1(rd_reg[59]), .A0N(N722), .A1N(n3850), .Y(
        N739) );
  OAI2BB2XL U593 ( .B0(n3690), .B1(rd_reg[58]), .A0N(N721), .A1N(n3850), .Y(
        N738) );
  OAI2BB2XL U594 ( .B0(n3700), .B1(rd_reg[57]), .A0N(N720), .A1N(n3850), .Y(
        N737) );
  OAI2BB2XL U595 ( .B0(n3700), .B1(rd_reg[56]), .A0N(N719), .A1N(n3850), .Y(
        N736) );
  OAI2BB2XL U596 ( .B0(n3670), .B1(rd_reg[45]), .A0N(N774), .A1N(n3760), .Y(
        N791) );
  OAI2BB2XL U597 ( .B0(n3680), .B1(rd_reg[44]), .A0N(N773), .A1N(n3750), .Y(
        N790) );
  OAI2BB2XL U598 ( .B0(n3670), .B1(rd_reg[43]), .A0N(N772), .A1N(n3760), .Y(
        N789) );
  OAI2BB2XL U599 ( .B0(n3670), .B1(rd_reg[42]), .A0N(N771), .A1N(n3750), .Y(
        N788) );
  OAI2BB2XL U600 ( .B0(n3670), .B1(rd_reg[41]), .A0N(N770), .A1N(n3870), .Y(
        N787) );
  OAI2BB2XL U601 ( .B0(n3670), .B1(rd_reg[40]), .A0N(N769), .A1N(n3870), .Y(
        N786) );
  OAI2BB2XL U602 ( .B0(n3700), .B1(rd_reg[28]), .A0N(N823), .A1N(n3790), .Y(
        N840) );
  OAI2BB2XL U603 ( .B0(n3700), .B1(rd_reg[27]), .A0N(N822), .A1N(n3780), .Y(
        N839) );
  OAI2BB2XL U604 ( .B0(n3700), .B1(rd_reg[26]), .A0N(N821), .A1N(n3780), .Y(
        N838) );
  OAI2BB2XL U605 ( .B0(n3690), .B1(rd_reg[25]), .A0N(N820), .A1N(n3780), .Y(
        N837) );
  OAI2BB2XL U606 ( .B0(n3690), .B1(rd_reg[24]), .A0N(N819), .A1N(n3780), .Y(
        N836) );
  OAI2BB2XL U607 ( .B0(n12), .B1(n345), .A0N(N56), .A1N(n345), .Y(n1083) );
  ADDHXL U608 ( .A(N9040), .B(N9030), .CO(add_101_aco_carry[2]), .S(N40) );
  ADDHXL U609 ( .A(N9050), .B(add_101_aco_carry[2]), .CO(add_101_aco_carry[3]), 
        .S(N41) );
  AO22X1 U610 ( .A0(n1930), .A1(rd_addr[9]), .B0(N57), .B1(n346), .Y(n1082) );
  ADDHXL U611 ( .A(N9060), .B(add_101_aco_carry[3]), .CO(add_101_aco_carry[4]), 
        .S(N42) );
  OAI21X1 U612 ( .A0(cnt[4]), .A1(n1930), .B0(n2810), .Y(n2740) );
  NAND3X1 U613 ( .A(out_cs[1]), .B(n86), .C(Vsync), .Y(n2810) );
  NOR2BX1 U614 ( .AN(n2800), .B(n2740), .Y(n2750) );
  OAI22XL U615 ( .A0(n4840), .A1(n700), .B0(n451), .B1(n701), .Y(n941) );
  OAI22XL U616 ( .A0(n4860), .A1(n8110), .B0(n4600), .B1(n8270), .Y(n8130) );
  OAI22XL U617 ( .A0(n4880), .A1(n800), .B0(n4610), .B1(n801), .Y(n8240) );
  OAI22XL U618 ( .A0(n4880), .A1(n798), .B0(n4610), .B1(n799), .Y(n8290) );
  OAI22XL U619 ( .A0(n4890), .A1(n7840), .B0(n4620), .B1(n7850), .Y(n845) );
  OAI22XL U620 ( .A0(n4910), .A1(n7700), .B0(n4630), .B1(n7710), .Y(n8610) );
  OAI22XL U621 ( .A0(n4920), .A1(n756), .B0(n4650), .B1(n757), .Y(n8770) );
  OAI22XL U622 ( .A0(n495), .A1(n7420), .B0(n4660), .B1(n7430), .Y(n8930) );
  OAI22XL U623 ( .A0(n4840), .A1(n98), .B0(n452), .B1(n702), .Y(n938) );
  OAI22XL U624 ( .A0(n4770), .A1(n99), .B0(n452), .B1(n6880), .Y(n954) );
  OAI22XL U625 ( .A0(n4770), .A1(n6860), .B0(n453), .B1(n6870), .Y(n957) );
  OAI22XL U626 ( .A0(n4780), .A1(n100), .B0(n454), .B1(n6740), .Y(n970) );
  OAI22XL U627 ( .A0(n4780), .A1(n6720), .B0(n454), .B1(n6730), .Y(n973) );
  OAI22XL U628 ( .A0(n4800), .A1(n101), .B0(n455), .B1(n6600), .Y(n986) );
  OAI22XL U629 ( .A0(n4800), .A1(n658), .B0(n455), .B1(n659), .Y(n989) );
  OAI22XL U630 ( .A0(n4810), .A1(n102), .B0(n456), .B1(n646), .Y(n1002) );
  OAI22XL U631 ( .A0(n4810), .A1(n644), .B0(n456), .B1(n645), .Y(n1005) );
  OAI22XL U632 ( .A0(n4830), .A1(n103), .B0(n457), .B1(n6320), .Y(n1018) );
  OAI22XL U633 ( .A0(n4830), .A1(n6300), .B0(n457), .B1(n6310), .Y(n1021) );
  OAI22XL U634 ( .A0(n4840), .A1(n97), .B0(n458), .B1(n6180), .Y(n1034) );
  OAI22XL U635 ( .A0(n4840), .A1(n6160), .B0(n458), .B1(n6170), .Y(n1037) );
  OAI22XL U636 ( .A0(n4850), .A1(n105), .B0(n459), .B1(n604), .Y(n1050) );
  OAI22XL U637 ( .A0(n4850), .A1(n602), .B0(n459), .B1(n603), .Y(n1053) );
  OAI22XL U638 ( .A0(n507), .A1(n7280), .B0(n4670), .B1(n7290), .Y(n909) );
  OAI22XL U639 ( .A0(n497), .A1(n104), .B0(n4670), .B1(n7160), .Y(n922) );
  OAI22XL U640 ( .A0(n497), .A1(n7140), .B0(n4680), .B1(n7150), .Y(n925) );
  NOR3X1 U641 ( .A(n86), .B(out_cs[2]), .C(n88), .Y(n1075) );
  OAI2BB2XL U642 ( .B0(n8), .B1(n345), .A0N(N52), .A1N(n345), .Y(n1087) );
  OAI2BB2XL U643 ( .B0(n3720), .B1(rd_reg[8]), .A0N(N868), .A1N(n3790), .Y(
        N885) );
  OAI2BB2XL U644 ( .B0(n3720), .B1(rd_reg[7]), .A0N(N867), .A1N(n3790), .Y(
        N884) );
  OAI2BB2XL U645 ( .B0(n3720), .B1(rd_reg[6]), .A0N(N866), .A1N(n3800), .Y(
        N883) );
  OAI2BB2XL U646 ( .B0(n3650), .B1(rd_reg[231]), .A0N(N168), .A1N(n3800), .Y(
        N185) );
  OAI2BB2XL U647 ( .B0(n3650), .B1(rd_reg[230]), .A0N(N167), .A1N(n3800), .Y(
        N184) );
  OAI2BB2XL U648 ( .B0(n3650), .B1(rd_reg[229]), .A0N(N166), .A1N(n3800), .Y(
        N183) );
  OAI2BB2XL U649 ( .B0(n3650), .B1(rd_reg[228]), .A0N(N165), .A1N(n3800), .Y(
        N182) );
  OAI2BB2XL U650 ( .B0(n3650), .B1(rd_reg[227]), .A0N(N164), .A1N(n3750), .Y(
        N181) );
  OAI2BB2XL U651 ( .B0(n3650), .B1(rd_reg[226]), .A0N(N163), .A1N(n3800), .Y(
        N180) );
  OAI2BB2XL U652 ( .B0(n3650), .B1(rd_reg[225]), .A0N(N162), .A1N(n3800), .Y(
        N179) );
  OAI2BB2XL U653 ( .B0(n3660), .B1(rd_reg[224]), .A0N(N161), .A1N(n3800), .Y(
        N178) );
  OAI2BB2XL U654 ( .B0(n3660), .B1(rd_reg[223]), .A0N(N160), .A1N(n3790), .Y(
        N177) );
  OAI2BB2XL U655 ( .B0(n3690), .B1(rd_reg[31]), .A0N(N760), .A1N(n3860), .Y(
        N777) );
  OAI2BB2XL U656 ( .B0(n3710), .B1(rd_reg[0]), .A0N(N860), .A1N(n3790), .Y(
        N877) );
  OAI2BB2XL U657 ( .B0(n3670), .B1(rd_reg[15]), .A0N(N810), .A1N(n3760), .Y(
        N827) );
  OAI2BB2XL U658 ( .B0(n3740), .B1(rd_reg[66]), .A0N(N663), .A1N(n3810), .Y(
        N680) );
  OAI2BB2XL U659 ( .B0(n3740), .B1(rd_reg[65]), .A0N(N662), .A1N(n3810), .Y(
        N679) );
  OAI2BB2XL U660 ( .B0(n3660), .B1(rd_reg[247]), .A0N(N118), .A1N(n3770), .Y(
        N135) );
  OAI2BB2XL U661 ( .B0(n3660), .B1(rd_reg[246]), .A0N(N117), .A1N(n3770), .Y(
        N134) );
  OAI2BB2XL U662 ( .B0(n3660), .B1(rd_reg[245]), .A0N(N116), .A1N(n3760), .Y(
        N133) );
  OAI2BB2XL U663 ( .B0(n3670), .B1(rd_reg[244]), .A0N(N115), .A1N(n3760), .Y(
        N132) );
  OAI2BB2XL U664 ( .B0(n3670), .B1(rd_reg[243]), .A0N(N114), .A1N(n3760), .Y(
        N131) );
  OAI2BB2XL U665 ( .B0(n3670), .B1(rd_reg[242]), .A0N(N113), .A1N(n3760), .Y(
        N130) );
  OAI2BB2XL U666 ( .B0(n3670), .B1(rd_reg[241]), .A0N(N112), .A1N(n3750), .Y(
        N129) );
  OAI2BB2XL U667 ( .B0(n353), .B1(rd_reg[240]), .A0N(N111), .A1N(n3760), .Y(
        N128) );
  OAI2BB2XL U668 ( .B0(n356), .B1(rd_reg[239]), .A0N(N110), .A1N(n3750), .Y(
        N127) );
  OAI2BB2XL U669 ( .B0(n3640), .B1(rd_reg[215]), .A0N(N218), .A1N(n3780), .Y(
        N235) );
  OAI2BB2XL U670 ( .B0(n3640), .B1(rd_reg[214]), .A0N(N217), .A1N(n3780), .Y(
        N234) );
  OAI2BB2XL U671 ( .B0(n3640), .B1(rd_reg[213]), .A0N(N216), .A1N(n3790), .Y(
        N233) );
  OAI2BB2XL U672 ( .B0(n3640), .B1(rd_reg[212]), .A0N(N215), .A1N(n3790), .Y(
        N232) );
  OAI2BB2XL U673 ( .B0(n3640), .B1(rd_reg[211]), .A0N(N214), .A1N(n3790), .Y(
        N231) );
  OAI2BB2XL U674 ( .B0(n3640), .B1(rd_reg[210]), .A0N(N213), .A1N(n3790), .Y(
        N230) );
  OAI2BB2XL U675 ( .B0(n3640), .B1(rd_reg[209]), .A0N(N212), .A1N(n3790), .Y(
        N229) );
  OAI2BB2XL U676 ( .B0(n3640), .B1(rd_reg[208]), .A0N(N211), .A1N(n3790), .Y(
        N228) );
  OAI2BB2XL U677 ( .B0(n3640), .B1(rd_reg[207]), .A0N(N210), .A1N(n3790), .Y(
        N227) );
  OAI2BB2XL U678 ( .B0(n3620), .B1(rd_reg[199]), .A0N(N268), .A1N(n3760), .Y(
        N285) );
  OAI2BB2XL U679 ( .B0(n3620), .B1(rd_reg[198]), .A0N(N267), .A1N(n3770), .Y(
        N284) );
  OAI2BB2XL U680 ( .B0(n3620), .B1(rd_reg[197]), .A0N(N266), .A1N(n3770), .Y(
        N283) );
  OAI2BB2XL U681 ( .B0(n3630), .B1(rd_reg[196]), .A0N(N265), .A1N(n3770), .Y(
        N282) );
  OAI2BB2XL U682 ( .B0(n3630), .B1(rd_reg[195]), .A0N(N264), .A1N(n3770), .Y(
        N281) );
  OAI2BB2XL U683 ( .B0(n3630), .B1(rd_reg[194]), .A0N(N263), .A1N(n3770), .Y(
        N280) );
  OAI2BB2XL U684 ( .B0(n3630), .B1(rd_reg[193]), .A0N(N262), .A1N(n3770), .Y(
        N279) );
  OAI2BB2XL U685 ( .B0(n3630), .B1(rd_reg[192]), .A0N(N261), .A1N(n3770), .Y(
        N278) );
  OAI2BB2XL U686 ( .B0(n3630), .B1(rd_reg[191]), .A0N(N260), .A1N(n3770), .Y(
        N277) );
  OAI2BB2XL U687 ( .B0(n3610), .B1(rd_reg[183]), .A0N(N318), .A1N(n3750), .Y(
        N335) );
  OAI2BB2XL U688 ( .B0(n3610), .B1(rd_reg[182]), .A0N(N317), .A1N(n3760), .Y(
        N334) );
  OAI2BB2XL U689 ( .B0(n3610), .B1(rd_reg[181]), .A0N(N316), .A1N(n3750), .Y(
        N333) );
  OAI2BB2XL U690 ( .B0(n3610), .B1(rd_reg[180]), .A0N(N315), .A1N(n3750), .Y(
        N332) );
  OAI2BB2XL U691 ( .B0(n3610), .B1(rd_reg[179]), .A0N(N314), .A1N(n3750), .Y(
        N331) );
  OAI2BB2XL U692 ( .B0(n3610), .B1(rd_reg[178]), .A0N(N313), .A1N(n3760), .Y(
        N330) );
  OAI2BB2XL U693 ( .B0(n3610), .B1(rd_reg[177]), .A0N(N312), .A1N(n3750), .Y(
        N329) );
  OAI2BB2XL U694 ( .B0(n3620), .B1(rd_reg[176]), .A0N(N311), .A1N(n3750), .Y(
        N328) );
  OAI2BB2XL U695 ( .B0(n3620), .B1(rd_reg[175]), .A0N(N310), .A1N(n3750), .Y(
        N327) );
  OAI2BB2XL U696 ( .B0(n3600), .B1(rd_reg[167]), .A0N(N368), .A1N(n3870), .Y(
        N385) );
  OAI2BB2XL U697 ( .B0(n3600), .B1(rd_reg[166]), .A0N(N367), .A1N(n3870), .Y(
        N384) );
  OAI2BB2XL U698 ( .B0(n3600), .B1(rd_reg[165]), .A0N(N366), .A1N(n3870), .Y(
        N383) );
  OAI2BB2XL U699 ( .B0(n3600), .B1(rd_reg[164]), .A0N(N365), .A1N(n3870), .Y(
        N382) );
  OAI2BB2XL U700 ( .B0(n3600), .B1(rd_reg[163]), .A0N(N364), .A1N(n3870), .Y(
        N381) );
  OAI2BB2XL U701 ( .B0(n3600), .B1(rd_reg[162]), .A0N(N363), .A1N(n3870), .Y(
        N380) );
  OAI2BB2XL U702 ( .B0(n3600), .B1(rd_reg[161]), .A0N(N362), .A1N(n3870), .Y(
        N379) );
  OAI2BB2XL U703 ( .B0(n3600), .B1(rd_reg[160]), .A0N(N361), .A1N(n3870), .Y(
        N378) );
  OAI2BB2XL U704 ( .B0(n3600), .B1(rd_reg[159]), .A0N(N360), .A1N(n3870), .Y(
        N377) );
  OAI2BB2XL U705 ( .B0(n358), .B1(rd_reg[151]), .A0N(N418), .A1N(n3850), .Y(
        N435) );
  OAI2BB2XL U706 ( .B0(n358), .B1(rd_reg[150]), .A0N(N417), .A1N(n3850), .Y(
        N434) );
  OAI2BB2XL U707 ( .B0(n358), .B1(rd_reg[149]), .A0N(N416), .A1N(n3850), .Y(
        N433) );
  OAI2BB2XL U708 ( .B0(n358), .B1(rd_reg[148]), .A0N(N415), .A1N(n3860), .Y(
        N432) );
  OAI2BB2XL U709 ( .B0(n359), .B1(rd_reg[147]), .A0N(N414), .A1N(n3860), .Y(
        N431) );
  OAI2BB2XL U710 ( .B0(n359), .B1(rd_reg[146]), .A0N(N413), .A1N(n3860), .Y(
        N430) );
  OAI2BB2XL U711 ( .B0(n359), .B1(rd_reg[145]), .A0N(N412), .A1N(n3860), .Y(
        N429) );
  OAI2BB2XL U712 ( .B0(n359), .B1(rd_reg[144]), .A0N(N411), .A1N(n3860), .Y(
        N428) );
  OAI2BB2XL U713 ( .B0(n359), .B1(rd_reg[143]), .A0N(N410), .A1N(n3860), .Y(
        N427) );
  OAI2BB2XL U714 ( .B0(n357), .B1(rd_reg[135]), .A0N(N468), .A1N(n3840), .Y(
        N485) );
  OAI2BB2XL U715 ( .B0(n357), .B1(rd_reg[134]), .A0N(N467), .A1N(n3840), .Y(
        N484) );
  OAI2BB2XL U716 ( .B0(n357), .B1(rd_reg[133]), .A0N(N466), .A1N(n3840), .Y(
        N483) );
  OAI2BB2XL U717 ( .B0(n357), .B1(rd_reg[132]), .A0N(N465), .A1N(n3840), .Y(
        N482) );
  OAI2BB2XL U718 ( .B0(n357), .B1(rd_reg[131]), .A0N(N464), .A1N(n3840), .Y(
        N481) );
  OAI2BB2XL U719 ( .B0(n357), .B1(rd_reg[130]), .A0N(N463), .A1N(n3850), .Y(
        N480) );
  OAI2BB2XL U720 ( .B0(n357), .B1(rd_reg[129]), .A0N(N462), .A1N(n3850), .Y(
        N479) );
  OAI2BB2XL U721 ( .B0(n357), .B1(rd_reg[128]), .A0N(N461), .A1N(n3850), .Y(
        N478) );
  OAI2BB2XL U722 ( .B0(n358), .B1(rd_reg[127]), .A0N(N460), .A1N(n3850), .Y(
        N477) );
  OAI2BB2XL U723 ( .B0(n356), .B1(rd_reg[119]), .A0N(N518), .A1N(n3830), .Y(
        N535) );
  OAI2BB2XL U724 ( .B0(n356), .B1(rd_reg[118]), .A0N(N517), .A1N(n3830), .Y(
        N534) );
  OAI2BB2XL U725 ( .B0(n356), .B1(rd_reg[117]), .A0N(N516), .A1N(n3830), .Y(
        N533) );
  OAI2BB2XL U726 ( .B0(n356), .B1(rd_reg[116]), .A0N(N515), .A1N(n3830), .Y(
        N532) );
  OAI2BB2XL U727 ( .B0(n356), .B1(rd_reg[115]), .A0N(N514), .A1N(n3830), .Y(
        N531) );
  OAI2BB2XL U728 ( .B0(n356), .B1(rd_reg[114]), .A0N(N513), .A1N(n3830), .Y(
        N530) );
  OAI2BB2XL U729 ( .B0(n356), .B1(rd_reg[113]), .A0N(N512), .A1N(n3830), .Y(
        N529) );
  OAI2BB2XL U730 ( .B0(n356), .B1(rd_reg[112]), .A0N(N511), .A1N(n3800), .Y(
        N528) );
  OAI2BB2XL U731 ( .B0(n3670), .B1(rd_reg[111]), .A0N(N510), .A1N(n3830), .Y(
        N527) );
  OAI2BB2XL U732 ( .B0(n354), .B1(rd_reg[103]), .A0N(N568), .A1N(n3820), .Y(
        N585) );
  OAI2BB2XL U733 ( .B0(n354), .B1(rd_reg[102]), .A0N(N567), .A1N(n3820), .Y(
        N584) );
  OAI2BB2XL U734 ( .B0(n354), .B1(rd_reg[101]), .A0N(N566), .A1N(n3820), .Y(
        N583) );
  OAI2BB2XL U735 ( .B0(n354), .B1(rd_reg[100]), .A0N(N565), .A1N(n3820), .Y(
        N582) );
  OAI2BB2XL U736 ( .B0(n355), .B1(rd_reg[99]), .A0N(N564), .A1N(n3820), .Y(
        N581) );
  OAI2BB2XL U737 ( .B0(n355), .B1(rd_reg[98]), .A0N(N563), .A1N(n3820), .Y(
        N580) );
  OAI2BB2XL U738 ( .B0(n355), .B1(rd_reg[97]), .A0N(N562), .A1N(n3820), .Y(
        N579) );
  OAI2BB2XL U739 ( .B0(n355), .B1(rd_reg[96]), .A0N(N561), .A1N(n3820), .Y(
        N578) );
  OAI2BB2XL U740 ( .B0(n355), .B1(rd_reg[95]), .A0N(N560), .A1N(n3820), .Y(
        N577) );
  OAI2BB2XL U741 ( .B0(n353), .B1(rd_reg[87]), .A0N(N618), .A1N(n3810), .Y(
        N635) );
  OAI2BB2XL U742 ( .B0(n353), .B1(rd_reg[86]), .A0N(N617), .A1N(n3810), .Y(
        N634) );
  OAI2BB2XL U743 ( .B0(n353), .B1(rd_reg[85]), .A0N(N616), .A1N(n3810), .Y(
        N633) );
  OAI2BB2XL U744 ( .B0(n353), .B1(rd_reg[84]), .A0N(N615), .A1N(n3810), .Y(
        N632) );
  OAI2BB2XL U745 ( .B0(n353), .B1(rd_reg[83]), .A0N(N614), .A1N(n3810), .Y(
        N631) );
  OAI2BB2XL U746 ( .B0(n353), .B1(rd_reg[82]), .A0N(N613), .A1N(n3810), .Y(
        N630) );
  OAI2BB2XL U747 ( .B0(n353), .B1(rd_reg[81]), .A0N(N612), .A1N(n3810), .Y(
        N629) );
  OAI2BB2XL U748 ( .B0(n353), .B1(rd_reg[80]), .A0N(N611), .A1N(n3810), .Y(
        N628) );
  OAI2BB2XL U749 ( .B0(n354), .B1(rd_reg[79]), .A0N(N610), .A1N(n3810), .Y(
        N627) );
  OAI2BB2XL U750 ( .B0(n3730), .B1(rd_reg[71]), .A0N(N668), .A1N(n3820), .Y(
        N685) );
  OAI2BB2XL U751 ( .B0(n3730), .B1(rd_reg[70]), .A0N(N667), .A1N(n3820), .Y(
        N684) );
  OAI2BB2XL U752 ( .B0(n3730), .B1(rd_reg[69]), .A0N(N666), .A1N(n3820), .Y(
        N683) );
  OAI2BB2XL U753 ( .B0(n3730), .B1(rd_reg[68]), .A0N(N665), .A1N(n3820), .Y(
        N682) );
  OAI2BB2XL U754 ( .B0(n3730), .B1(rd_reg[67]), .A0N(N664), .A1N(n3820), .Y(
        N681) );
  OAI2BB2XL U755 ( .B0(n3730), .B1(rd_reg[64]), .A0N(N661), .A1N(n3810), .Y(
        N678) );
  OAI2BB2XL U756 ( .B0(n3730), .B1(rd_reg[63]), .A0N(N660), .A1N(n3810), .Y(
        N677) );
  OAI2BB2XL U757 ( .B0(n3700), .B1(rd_reg[55]), .A0N(N718), .A1N(n3850), .Y(
        N735) );
  OAI2BB2XL U758 ( .B0(n3700), .B1(rd_reg[54]), .A0N(N717), .A1N(n3840), .Y(
        N734) );
  OAI2BB2XL U759 ( .B0(n3700), .B1(rd_reg[53]), .A0N(N716), .A1N(n3840), .Y(
        N733) );
  OAI2BB2XL U760 ( .B0(n3700), .B1(rd_reg[52]), .A0N(N715), .A1N(n3840), .Y(
        N732) );
  OAI2BB2XL U761 ( .B0(n3700), .B1(rd_reg[51]), .A0N(N714), .A1N(n3840), .Y(
        N731) );
  OAI2BB2XL U762 ( .B0(n3710), .B1(rd_reg[50]), .A0N(N713), .A1N(n3840), .Y(
        N730) );
  OAI2BB2XL U763 ( .B0(n3710), .B1(rd_reg[49]), .A0N(N712), .A1N(n3840), .Y(
        N729) );
  OAI2BB2XL U764 ( .B0(n3710), .B1(rd_reg[48]), .A0N(N711), .A1N(n3840), .Y(
        N728) );
  OAI2BB2XL U765 ( .B0(n3710), .B1(rd_reg[47]), .A0N(N710), .A1N(n3830), .Y(
        N727) );
  OAI2BB2XL U766 ( .B0(n3680), .B1(rd_reg[39]), .A0N(N768), .A1N(n3870), .Y(
        N785) );
  OAI2BB2XL U767 ( .B0(n3680), .B1(rd_reg[38]), .A0N(N767), .A1N(n3870), .Y(
        N784) );
  OAI2BB2XL U768 ( .B0(n3680), .B1(rd_reg[37]), .A0N(N766), .A1N(n3870), .Y(
        N783) );
  OAI2BB2XL U769 ( .B0(n3680), .B1(rd_reg[36]), .A0N(N765), .A1N(n3870), .Y(
        N782) );
  OAI2BB2XL U770 ( .B0(n3680), .B1(rd_reg[35]), .A0N(N764), .A1N(n3860), .Y(
        N781) );
  OAI2BB2XL U771 ( .B0(n3680), .B1(rd_reg[34]), .A0N(N763), .A1N(n3860), .Y(
        N780) );
  OAI2BB2XL U772 ( .B0(n3680), .B1(rd_reg[33]), .A0N(N762), .A1N(n3860), .Y(
        N779) );
  OAI2BB2XL U773 ( .B0(n3690), .B1(rd_reg[32]), .A0N(N761), .A1N(n3860), .Y(
        N778) );
  OAI2BB2XL U774 ( .B0(n3690), .B1(rd_reg[23]), .A0N(N818), .A1N(n3780), .Y(
        N835) );
  OAI2BB2XL U775 ( .B0(n3690), .B1(rd_reg[22]), .A0N(N817), .A1N(n3770), .Y(
        N834) );
  OAI2BB2XL U776 ( .B0(n3690), .B1(rd_reg[21]), .A0N(N816), .A1N(n3770), .Y(
        N833) );
  OAI2BB2XL U777 ( .B0(n3680), .B1(rd_reg[20]), .A0N(N815), .A1N(n3770), .Y(
        N832) );
  OAI2BB2XL U778 ( .B0(n3680), .B1(rd_reg[19]), .A0N(N814), .A1N(n3770), .Y(
        N831) );
  OAI2BB2XL U779 ( .B0(n3680), .B1(rd_reg[18]), .A0N(N813), .A1N(n3760), .Y(
        N830) );
  OAI2BB2XL U780 ( .B0(n3680), .B1(rd_reg[17]), .A0N(N812), .A1N(n3760), .Y(
        N829) );
  OAI2BB2XL U781 ( .B0(n3720), .B1(rd_reg[16]), .A0N(N811), .A1N(n3760), .Y(
        N828) );
  OAI2BB2XL U782 ( .B0(n3720), .B1(rd_reg[5]), .A0N(N865), .A1N(n3800), .Y(
        N882) );
  OAI2BB2XL U783 ( .B0(n3710), .B1(rd_reg[4]), .A0N(N864), .A1N(n3800), .Y(
        N881) );
  OAI2BB2XL U784 ( .B0(n3710), .B1(rd_reg[3]), .A0N(N863), .A1N(n3800), .Y(
        N880) );
  OAI2BB2XL U785 ( .B0(n3710), .B1(rd_reg[2]), .A0N(N862), .A1N(n3800), .Y(
        N879) );
  OAI2BB2XL U786 ( .B0(n3710), .B1(rd_reg[1]), .A0N(N861), .A1N(n3800), .Y(
        N878) );
  OAI21XL U787 ( .A0(n2750), .A1(n96), .B0(n5870), .Y(n1093) );
  OAI2BB2XL U788 ( .B0(n11), .B1(n345), .A0N(N55), .A1N(n345), .Y(n1084) );
  OAI2BB2XL U789 ( .B0(n10), .B1(n346), .A0N(N54), .A1N(n346), .Y(n1085) );
  OAI2BB2XL U790 ( .B0(n9), .B1(n346), .A0N(N53), .A1N(n346), .Y(n1086) );
  OAI2BB2XL U791 ( .B0(n7), .B1(n345), .A0N(N51), .A1N(n345), .Y(n1088) );
  OAI2BB2XL U792 ( .B0(n6), .B1(n346), .A0N(N50), .A1N(n346), .Y(n1089) );
  OAI2BB2XL U793 ( .B0(n5), .B1(n346), .A0N(N49), .A1N(n346), .Y(n1090) );
  OAI2BB2XL U794 ( .B0(n4), .B1(n345), .A0N(N48), .A1N(n345), .Y(n1091) );
  OR3X2 U795 ( .A(out_cs[1]), .B(out_cs[2]), .C(n86), .Y(n1930) );
  AO22X1 U796 ( .A0(n4690), .A1(rd_reg[223]), .B0(n498), .B1(rd_reg[239]), .Y(
        n8120) );
  AO22X1 U797 ( .A0(n4690), .A1(rd_reg[227]), .B0(n498), .B1(rd_reg[243]), .Y(
        n8760) );
  AO22X1 U798 ( .A0(n4690), .A1(rd_reg[228]), .B0(n498), .B1(rd_reg[244]), .Y(
        n8920) );
  AO22X1 U799 ( .A0(n4690), .A1(rd_reg[230]), .B0(n498), .B1(rd_reg[246]), .Y(
        n924) );
  AO22X1 U800 ( .A0(n4690), .A1(rd_reg[231]), .B0(n498), .B1(rd_reg[247]), .Y(
        n940) );
  AO22X1 U801 ( .A0(n4690), .A1(rd_reg[232]), .B0(n498), .B1(rd_reg[248]), .Y(
        n956) );
  AO22X1 U802 ( .A0(n4690), .A1(rd_reg[236]), .B0(n498), .B1(rd_reg[252]), .Y(
        n1020) );
  AO22X1 U803 ( .A0(n4690), .A1(rd_reg[238]), .B0(n498), .B1(rd_reg[254]), .Y(
        n1052) );
  AO22X1 U804 ( .A0(n4690), .A1(rd_reg[226]), .B0(n497), .B1(rd_reg[242]), .Y(
        n8600) );
  AO22X1 U805 ( .A0(n4690), .A1(rd_reg[229]), .B0(n497), .B1(rd_reg[245]), .Y(
        n908) );
  AO22X1 U806 ( .A0(n4720), .A1(rd_reg[15]), .B0(n4690), .B1(rd_reg[0]), .Y(
        n8260) );
  AO22X1 U807 ( .A0(mode), .A1(rd_addr[10]), .B0(n5850), .B1(rd_addr[9]), .Y(
        N45) );
  CLKINVX1 U808 ( .A(mode), .Y(n5850) );
  AND2X1 U809 ( .A(cnt[0]), .B(Vsync), .Y(N9030) );
  AND2X1 U810 ( .A(cnt[1]), .B(Vsync), .Y(N9040) );
  AND2X1 U811 ( .A(cnt[2]), .B(Vsync), .Y(N9050) );
  AND2X1 U812 ( .A(cnt[3]), .B(Vsync), .Y(N9060) );
  AND2X1 U813 ( .A(Vsync), .B(cnt[4]), .Y(N9070) );
  CLKINVX1 U814 ( .A(N9030), .Y(N39) );
  XOR2X1 U815 ( .A(add_101_aco_carry[4]), .B(N9070), .Y(N43) );
  PWMConvert_DW01_inc_0 add_145_I16 ( .A({OUT[15], out_buffer[15:0]}), .SUM({
        N876, N875, N874, N873, N872, N871, N870, N869, N868, N867, N866, N865, 
        N864, N863, N862, N861, N860}) );
  PWMConvert_DW01_inc_1 add_145_I15 ( .A({OUT[14], out_buffer[31:16]}), .SUM({
        N826, N825, N824, N823, N822, N821, N820, N819, N818, N817, N816, N815, 
        N814, N813, N812, N811, N810}) );
  PWMConvert_DW01_inc_2 add_145_I14 ( .A({OUT[13], out_buffer[47:32]}), .SUM({
        N776, N775, N774, N773, N772, N771, N770, N769, N768, N767, N766, N765, 
        N764, N763, N762, N761, N760}) );
  PWMConvert_DW01_inc_3 add_145_I13 ( .A({OUT[12], out_buffer[63:48]}), .SUM({
        N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, 
        N714, N713, N712, N711, N710}) );
  PWMConvert_DW01_inc_4 add_145_I12 ( .A({OUT[11], out_buffer[79:64]}), .SUM({
        N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, N665, 
        N664, N663, N662, N661, N660}) );
  PWMConvert_DW01_inc_5 add_145_I11 ( .A({OUT[10], out_buffer[95:80]}), .SUM({
        N626, N625, N624, N623, N622, N621, N620, N619, N618, N617, N616, N615, 
        N614, N613, N612, N611, N610}) );
  PWMConvert_DW01_inc_6 add_145_I10 ( .A({OUT[9], out_buffer[111:96]}), .SUM({
        N576, N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, 
        N564, N563, N562, N561, N560}) );
  PWMConvert_DW01_inc_7 add_145_I9 ( .A({OUT[8], out_buffer[127:112]}), .SUM({
        N526, N525, N524, N523, N522, N521, N520, N519, N518, N517, N516, N515, 
        N514, N513, N512, N511, N510}) );
  PWMConvert_DW01_inc_8 add_145_I8 ( .A({OUT[7], out_buffer[143:128]}), .SUM({
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460}) );
  PWMConvert_DW01_inc_9 add_145_I7 ( .A({OUT[6], out_buffer[159:144]}), .SUM({
        N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, 
        N414, N413, N412, N411, N410}) );
  PWMConvert_DW01_inc_10 add_145_I6 ( .A({OUT[5], out_buffer[175:160]}), .SUM(
        {N376, N375, N374, N373, N372, N371, N370, N369, N368, N367, N366, 
        N365, N364, N363, N362, N361, N360}) );
  PWMConvert_DW01_inc_11 add_145_I5 ( .A({OUT[4], out_buffer[191:176]}), .SUM(
        {N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316, 
        N315, N314, N313, N312, N311, N310}) );
  PWMConvert_DW01_inc_12 add_145_I4 ( .A({OUT[3], out_buffer[207:192]}), .SUM(
        {N276, N275, N274, N273, N272, N271, N270, N269, N268, N267, N266, 
        N265, N264, N263, N262, N261, N260}) );
  PWMConvert_DW01_inc_13 add_145_I3 ( .A({OUT[2], out_buffer[223:208]}), .SUM(
        {N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, 
        N215, N214, N213, N212, N211, N210}) );
  PWMConvert_DW01_inc_14 add_145_I2 ( .A({OUT[1], out_buffer[239:224]}), .SUM(
        {N176, N175, N174, N173, N172, N171, N170, N169, N168, N167, N166, 
        N165, N164, N163, N162, N161, N160}) );
  PWMConvert_DW01_inc_15 add_145 ( .A({OUT[0], out_buffer[255:240]}), .SUM({
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110}) );
  PWMConvert_DW01_inc_16 add_116_S2 ( .A({rd_addr, addr}), .SUM({N58, N57, N56, 
        N55, N54, N53, N52, N51, N50, N49, N48}) );
endmodule


module LEDDC ( DCK, DAI, DEN, GCK, Vsync, mode, rst, OUT );
  output [15:0] OUT;
  input DCK, DAI, DEN, GCK, Vsync, mode, rst;
  wire   en_rd, en_wd1, en_wd2, n_1_net_, n4, n5, n6, n7, n8;
  wire   [15:0] rd_data;
  wire   [15:0] rd_data1;
  wire   [15:0] rd_data2;
  wire   [8:0] wd_addr;
  wire   [15:0] r_data;
  wire   [8:0] rd_addr;

  sram_512x16 ram1 ( .AB(wd_addr), .DB(r_data), .AA(rd_addr), .QA(rd_data1), 
        .CENB(en_wd1), .CENA(n5), .CLKB(n_1_net_), .CLKA(GCK) );
  sram_512x16 ram2 ( .AB(wd_addr), .DB(r_data), .AA(rd_addr), .QA(rd_data2), 
        .CENB(en_wd2), .CENA(n8), .CLKB(n_1_net_), .CLKA(GCK) );
  CLKINVX6 U17 ( .A(DCK), .Y(n_1_net_) );
  NAND2X4 U19 ( .A(n6), .B(n7), .Y(rd_data[3]) );
  NAND2X2 U20 ( .A(rd_data2[3]), .B(n5), .Y(n6) );
  NAND2X2 U21 ( .A(rd_data1[3]), .B(n8), .Y(n7) );
  CLKMX2X2 U22 ( .A(rd_data2[4]), .B(rd_data1[4]), .S0(n8), .Y(rd_data[4]) );
  CLKMX2X2 U23 ( .A(rd_data2[8]), .B(rd_data1[8]), .S0(n8), .Y(rd_data[8]) );
  CLKMX2X4 U24 ( .A(rd_data2[1]), .B(rd_data1[1]), .S0(n8), .Y(rd_data[1]) );
  CLKMX2X2 U25 ( .A(rd_data2[5]), .B(rd_data1[5]), .S0(n8), .Y(rd_data[5]) );
  BUFX4 U26 ( .A(en_rd), .Y(n8) );
  BUFX2 U27 ( .A(DAI), .Y(n4) );
  CLKMX2X6 U28 ( .A(rd_data2[0]), .B(rd_data1[0]), .S0(n8), .Y(rd_data[0]) );
  INVX1 U29 ( .A(n8), .Y(n5) );
  CLKMX2X2 U30 ( .A(rd_data2[10]), .B(rd_data1[10]), .S0(n8), .Y(rd_data[10])
         );
  MX2X1 U31 ( .A(rd_data2[11]), .B(rd_data1[11]), .S0(n8), .Y(rd_data[11]) );
  MX2X1 U32 ( .A(rd_data2[13]), .B(rd_data1[13]), .S0(n8), .Y(rd_data[13]) );
  MX2X1 U33 ( .A(rd_data2[12]), .B(rd_data1[12]), .S0(n8), .Y(rd_data[12]) );
  MX2XL U34 ( .A(rd_data2[14]), .B(rd_data1[14]), .S0(n8), .Y(rd_data[14]) );
  CLKMX2X2 U35 ( .A(rd_data2[7]), .B(rd_data1[7]), .S0(n8), .Y(rd_data[7]) );
  CLKMX2X2 U36 ( .A(rd_data2[6]), .B(rd_data1[6]), .S0(n8), .Y(rd_data[6]) );
  CLKMX2X2 U37 ( .A(rd_data2[9]), .B(rd_data1[9]), .S0(n8), .Y(rd_data[9]) );
  MX2XL U38 ( .A(rd_data2[15]), .B(rd_data1[15]), .S0(n8), .Y(rd_data[15]) );
  CLKMX2X2 U39 ( .A(rd_data2[2]), .B(rd_data1[2]), .S0(n8), .Y(rd_data[2]) );
  DataReceiver dr ( .DCK(DCK), .DAI(n4), .DEN(DEN), .rst(rst), .addr(wd_addr), 
        .data(r_data), .en1(en_wd1), .en2(en_wd2) );
  PWMConvert pc ( .GCK(GCK), .Vsync(Vsync), .mode(mode), .rst(rst), .OUT(OUT), 
        .data(rd_data), .addr(rd_addr), .en(en_rd) );
endmodule

